--
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes,",
--		 constants, and functions",
--

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package rom_pack is

  type RomType is array (natural range <>) of std_logic_vector(9 downto 0);

  constant ROM_35 : RomType := (
    8#0000# => '0' & O"335",
    8#0001# => '1' & O"377",
    8#0002# => '1' & O"044",
    8#0003# => '0' & O"027",
    8#0004# => '0' & O"504",
    8#0005# => '1' & O"104",
    8#0006# => '0' & O"204",
    8#0007# => '0' & O"420",
    8#0010# => '1' & O"321",
    8#0011# => '1' & O"773",
    8#0012# => '0' & O"137",
    8#0013# => '0' & O"303",
    8#0014# => '0' & O"650",
    8#0015# => '1' & O"547",
    8#0016# => '1' & O"356",
    8#0017# => '1' & O"742",
    8#0020# => '0' & O"056",
    8#0021# => '0' & O"220",
    8#0022# => '1' & O"752",
    8#0023# => '1' & O"752",
    8#0024# => '1' & O"752",
    8#0025# => '0' & O"153",
    8#0026# => '1' & O"151",
    8#0027# => '0' & O"250",
    8#0030# => '1' & O"250",
    8#0031# => '0' & O"377",
    8#0032# => '1' & O"752",
    8#0033# => '1' & O"752",
    8#0034# => '1' & O"752",
    8#0035# => '0' & O"060",
    8#0036# => '0' & O"314",
    8#0037# => '0' & O"252",
    8#0040# => '0' & O"650",
    8#0041# => '0' & O"103",
    8#0042# => '0' & O"723",
    8#0043# => '0' & O"314",
    8#0044# => '0' & O"060",
    8#0045# => '0' & O"000",
    8#0046# => '0' & O"203",
    8#0047# => '0' & O"504",
    8#0050# => '0' & O"104",
    8#0051# => '0' & O"273",
    8#0052# => '1' & O"104",
    8#0053# => '0' & O"237",
    8#0054# => '1' & O"204",
    8#0055# => '1' & O"413",
    8#0056# => '0' & O"056",
    8#0057# => '0' & O"220",
    8#0060# => '1' & O"450",
    8#0061# => '1' & O"557",
    8#0062# => '1' & O"752",
    8#0063# => '1' & O"752",
    8#0064# => '1' & O"752",
    8#0065# => '0' & O"113",
    8#0066# => '1' & O"147",
    8#0067# => '1' & O"650",
    8#0070# => '0' & O"561",
    8#0071# => '1' & O"567",
    8#0072# => '1' & O"713",
    8#0073# => '1' & O"316",
    8#0074# => '0' & O"304",
    8#0075# => '0' & O"733",
    8#0076# => '0' & O"450",
    8#0077# => '0' & O"064",
    8#0100# => '1' & O"316",
    8#0101# => '1' & O"565",
    8#0102# => '0' & O"456",
    8#0103# => '1' & O"372",
    8#0104# => '0' & O"426",
    8#0105# => '1' & O"552",
    8#0106# => '1' & O"603",
    8#0107# => '0' & O"672",
    8#0110# => '1' & O"633",
    8#0111# => '1' & O"466",
    8#0112# => '1' & O"514",
    8#0113# => '1' & O"633",
    8#0114# => '0' & O"034",
    8#0115# => '0' & O"752",
    8#0116# => '0' & O"002",
    8#0117# => '0' & O"463",
    8#0120# => '1' & O"304",
    8#0121# => '1' & O"326",
    8#0122# => '1' & O"646",
    8#0123# => '0' & O"424",
    8#0124# => '1' & O"037",
    8#0125# => '0' & O"575",
    8#0126# => '1' & O"567",
    8#0127# => '0' & O"322",
    8#0130# => '0' & O"562",
    8#0131# => '0' & O"332",
    8#0132# => '1' & O"612",
    8#0133# => '0' & O"567",
    8#0134# => '0' & O"316",
    8#0135# => '0' & O"064",
    8#0136# => '0' & O"616",
    8#0137# => '1' & O"414",
    8#0140# => '0' & O"452",
    8#0141# => '0' & O"612",
    8#0142# => '0' & O"672",
    8#0143# => '0' & O"643",
    8#0144# => '0' & O"252",
    8#0145# => '0' & O"572",
    8#0146# => '0' & O"537",
    8#0147# => '0' & O"514",
    8#0150# => '1' & O"652",
    8#0151# => '0' & O"424",
    8#0152# => '0' & O"413",
    8#0153# => '1' & O"452",
    8#0154# => '0' & O"052",
    8#0155# => '1' & O"735",
    8#0156# => '0' & O"412",
    8#0157# => '1' & O"316",
    8#0160# => '1' & O"454",
    8#0161# => '1' & O"047",
    8#0162# => '1' & O"662",
    8#0163# => '0' & O"753",
    8#0164# => '1' & O"321",
    8#0165# => '0' & O"220",
    8#0166# => '0' & O"424",
    8#0167# => '1' & O"733",
    8#0170# => '1' & O"662",
    8#0171# => '0' & O"372",
    8#0172# => '0' & O"616",
    8#0173# => '0' & O"672",
    8#0174# => '0' & O"777",
    8#0175# => '0' & O"332",
    8#0176# => '0' & O"252",
    8#0177# => '1' & O"514",
    8#0200# => '0' & O"426",
    8#0201# => '0' & O"552",
    8#0202# => '1' & O"176",
    8#0203# => '0' & O"473",
    8#0204# => '1' & O"166",
    8#0205# => '1' & O"003",
    8#0206# => '0' & O"312",
    8#0207# => '1' & O"735",
    8#0210# => '1' & O"326",
    8#0211# => '0' & O"636",
    8#0212# => '1' & O"454",
    8#0213# => '1' & O"117",
    8#0214# => '0' & O"216",
    8#0215# => '0' & O"756",
    8#0216# => '0' & O"114",
    8#0217# => '0' & O"422",
    8#0220# => '0' & O"074",
    8#0221# => '0' & O"642",
    8#0222# => '1' & O"077",
    8#0223# => '1' & O"656",
    8#0224# => '0' & O"354",
    8#0225# => '1' & O"747",
    8#0226# => '0' & O"312",
    8#0227# => '0' & O"604",
    8#0230# => '0' & O"753",
    8#0231# => '0' & O"376",
    8#0232# => '0' & O"650",
    8#0233# => '0' & O"056",
    8#0234# => '1' & O"772",
    8#0235# => '1' & O"772",
    8#0236# => '0' & O"772",
    8#0237# => '0' & O"772",
    8#0240# => '0' & O"112",
    8#0241# => '1' & O"217",
    8#0242# => '1' & O"656",
    8#0243# => '1' & O"646",
    8#0244# => '0' & O"646",
    8#0245# => '1' & O"237",
    8#0246# => '1' & O"656",
    8#0247# => '1' & O"046",
    8#0250# => '0' & O"112",
    8#0251# => '1' & O"373",
    8#0252# => '1' & O"216",
    8#0253# => '1' & O"752",
    8#0254# => '0' & O"016",
    8#0255# => '1' & O"373",
    8#0256# => '1' & O"243",
    8#0257# => '1' & O"366",
    8#0260# => '0' & O"324",
    8#0261# => '1' & O"323",
    8#0262# => '1' & O"576",
    8#0263# => '0' & O"376",
    8#0264# => '0' & O"724",
    8#0265# => '1' & O"337",
    8#0266# => '0' & O"450",
    8#0267# => '0' & O"704",
    8#0270# => '0' & O"316",
    8#0271# => '0' & O"556",
    8#0272# => '0' & O"276",
    8#0273# => '0' & O"776",
    8#0274# => '1' & O"056",
    8#0275# => '0' & O"060",
    8#0276# => '0' & O"220",
    8#0277# => '0' & O"561",
    8#0300# => '0' & O"504",
    8#0301# => '1' & O"567",
    8#0302# => '1' & O"316",
    8#0303# => '0' & O"636",
    8#0304# => '1' & O"044",
    8#0305# => '1' & O"477",
    8#0306# => '0' & O"772",
    8#0307# => '1' & O"004",
    8#0310# => '0' & O"524",
    8#0311# => '1' & O"467",
    8#0312# => '0' & O"752",
    8#0313# => '1' & O"433",
    8#0314# => '0' & O"050",
    8#0315# => '0' & O"024",
    8#0316# => '1' & O"437",
    8#0317# => '0' & O"044",
    8#0320# => '0' & O"034",
    8#0321# => '1' & O"454",
    8#0322# => '1' & O"503",
    8#0323# => '1' & O"050",
    8#0324# => '1' & O"024",
    8#0325# => '1' & O"463",
    8#0326# => '0' & O"416",
    8#0327# => '0' & O"544",
    8#0330# => '0' & O"320",
    8#0331# => '0' & O"450",
    8#0332# => '1' & O"656",
    8#0333# => '0' & O"565",
    8#0334# => '0' & O"704",
    8#0335# => '1' & O"735",
    8#0336# => '1' & O"275",
    8#0337# => '1' & O"053",
    8#0340# => '1' & O"326",
    8#0341# => '0' & O"034",
    8#0342# => '0' & O"254",
    8#0343# => '0' & O"427",
    8#0344# => '1' & O"414",
    8#0345# => '1' & O"356",
    8#0346# => '1' & O"366",
    8#0347# => '1' & O"742",
    8#0350# => '1' & O"742",
    8#0351# => '0' & O"214",
    8#0352# => '0' & O"074",
    8#0353# => '1' & O"542",
    8#0354# => '1' & O"677",
    8#0355# => '0' & O"002",
    8#0356# => '1' & O"653",
    8#0357# => '1' & O"742",
    8#0360# => '1' & O"456",
    8#0361# => '0' & O"060",
    8#0362# => '0' & O"404",
    8#0363# => '1' & O"324",
    8#0364# => '0' & O"163",
    8#0365# => '0' & O"677",
    8#0366# => '0' & O"376",
    8#0367# => '1' & O"244",
    8#0370# => '1' & O"417",
    8#0371# => '0' & O"624",
    8#0372# => '1' & O"763",
    8#0373# => '0' & O"034",
    8#0374# => '1' & O"222",
    8#0375# => '0' & O"751",
    8#0376# => '1' & O"250",
    8#0377# => '1' & O"557",
    8#0400# => '1' & O"717",
    8#0401# => '1' & O"456",
    8#0402# => '0' & O"241",
    8#0403# => '0' & O"650",
    8#0404# => '0' & O"241",
    8#0405# => '0' & O"650",
    8#0406# => '1' & O"124",
    8#0407# => '0' & O"047",
    8#0410# => '1' & O"656",
    8#0411# => '0' & O"524",
    8#0412# => '0' & O"113",
    8#0413# => '0' & O"336",
    8#0414# => '1' & O"231",
    8#0415# => '0' & O"450",
    8#0416# => '1' & O"225",
    8#0417# => '1' & O"141",
    8#0420# => '0' & O"225",
    8#0421# => '0' & O"650",
    8#0422# => '1' & O"231",
    8#0423# => '1' & O"224",
    8#0424# => '1' & O"553",
    8#0425# => '1' & O"356",
    8#0426# => '1' & O"742",
    8#0427# => '0' & O"446",
    8#0430# => '1' & O"646",
    8#0431# => '0' & O"552",
    8#0432# => '1' & O"222",
    8#0433# => '0' & O"672",
    8#0434# => '0' & O"147",
    8#0435# => '1' & O"322",
    8#0436# => '0' & O"752",
    8#0437# => '0' & O"167",
    8#0440# => '1' & O"316",
    8#0441# => '1' & O"216",
    8#0442# => '0' & O"450",
    8#0443# => '1' & O"056",
    8#0444# => '0' & O"407",
    8#0445# => '1' & O"056",
    8#0446# => '0' & O"414",
    8#0447# => '1' & O"573",
    8#0450# => '0' & O"450",
    8#0451# => '1' & O"656",
    8#0452# => '0' & O"642",
    8#0453# => '0' & O"267",
    8#0454# => '0' & O"256",
    8#0455# => '0' & O"616",
    8#0456# => '0' & O"212",
    8#0457# => '1' & O"457",
    8#0460# => '0' & O"616",
    8#0461# => '0' & O"124",
    8#0462# => '0' & O"227",
    8#0463# => '1' & O"224",
    8#0464# => '0' & O"667",
    8#0465# => '0' & O"524",
    8#0466# => '0' & O"127",
    8#0467# => '0' & O"376",
    8#0470# => '1' & O"676",
    8#0471# => '0' & O"067",
    8#0472# => '1' & O"222",
    8#0473# => '1' & O"576",
    8#0474# => '0' & O"353",
    8#0475# => '0' & O"776",
    8#0476# => '1' & O"462",
    8#0477# => '0' & O"722",
    8#0500# => '1' & O"456",
    8#0501# => '0' & O"456",
    8#0502# => '1' & O"522",
    8#0503# => '0' & O"357",
    8#0504# => '0' & O"650",
    8#0505# => '1' & O"316",
    8#0506# => '1' & O"662",
    8#0507# => '1' & O"456",
    8#0510# => '0' & O"422",
    8#0511# => '0' & O"450",
    8#0512# => '1' & O"776",
    8#0513# => '1' & O"776",
    8#0514# => '0' & O"217",
    8#0515# => '0' & O"316",
    8#0516# => '0' & O"052",
    8#0517# => '1' & O"326",
    8#0520# => '1' & O"311",
    8#0521# => '0' & O"542",
    8#0522# => '0' & O"650",
    8#0523# => '1' & O"656",
    8#0524# => '0' & O"414",
    8#0525# => '1' & O"221",
    8#0526# => '0' & O"614",
    8#0527# => '1' & O"155",
    8#0530# => '1' & O"014",
    8#0531# => '1' & O"155",
    8#0532# => '0' & O"214",
    8#0533# => '1' & O"030",
    8#0534# => '1' & O"214",
    8#0535# => '1' & O"155",
    8#0536# => '1' & O"071",
    8#0537# => '1' & O"155",
    8#0540# => '1' & O"461",
    8#0541# => '0' & O"416",
    8#0542# => '1' & O"155",
    8#0543# => '0' & O"216",
    8#0544# => '1' & O"455",
    8#0545# => '1' & O"461",
    8#0546# => '1' & O"256",
    8#0547# => '1' & O"231",
    8#0550# => '1' & O"124",
    8#0551# => '0' & O"663",
    8#0552# => '0' & O"376",
    8#0553# => '1' & O"141",
    8#0554# => '0' & O"144",
    8#0555# => '0' & O"316",
    8#0556# => '0' & O"542",
    8#0557# => '0' & O"752",
    8#0560# => '0' & O"124",
    8#0561# => '1' & O"227",
    8#0562# => '1' & O"231",
    8#0563# => '1' & O"461",
    8#0564# => '1' & O"256",
    8#0565# => '1' & O"225",
    8#0566# => '1' & O"461",
    8#0567# => '1' & O"256",
    8#0570# => '1' & O"256",
    8#0571# => '1' & O"125",
    8#0572# => '1' & O"256",
    8#0573# => '1' & O"655",
    8#0574# => '1' & O"461",
    8#0575# => '1' & O"214",
    8#0576# => '1' & O"161",
    8#0577# => '1' & O"071",
    8#0600# => '1' & O"014",
    8#0601# => '1' & O"165",
    8#0602# => '0' & O"214",
    8#0603# => '1' & O"030",
    8#0604# => '0' & O"614",
    8#0605# => '1' & O"161",
    8#0606# => '0' & O"414",
    8#0607# => '1' & O"161",
    8#0610# => '1' & O"161",
    8#0611# => '1' & O"456",
    8#0612# => '1' & O"116",
    8#0613# => '1' & O"514",
    8#0614# => '0' & O"530",
    8#0615# => '1' & O"757",
    8#0616# => '0' & O"614",
    8#0617# => '1' & O"030",
    8#0620# => '0' & O"630",
    8#0621# => '0' & O"530",
    8#0622# => '0' & O"230",
    8#0623# => '0' & O"430",
    8#0624# => '1' & O"130",
    8#0625# => '0' & O"124",
    8#0626# => '1' & O"553",
    8#0627# => '0' & O"060",
    8#0630# => '1' & O"356",
    8#0631# => '1' & O"742",
    8#0632# => '0' & O"020",
    8#0633# => '0' & O"420",
    8#0634# => '0' & O"416",
    8#0635# => '1' & O"226",
    8#0636# => '1' & O"056",
    8#0637# => '1' & O"207",
    8#0640# => '0' & O"776",
    8#0641# => '1' & O"416",
    8#0642# => '1' & O"203",
    8#0643# => '1' & O"616",
    8#0644# => '0' & O"420",
    8#0645# => '0' & O"420",
    8#0646# => '0' & O"512",
    8#0647# => '0' & O"420",
    8#0650# => '0' & O"742",
    8#0651# => '1' & O"516",
    8#0652# => '1' & O"243",
    8#0653# => '1' & O"716",
    8#0654# => '0' & O"416",
    8#0655# => '0' & O"034",
    8#0656# => '1' & O"122",
    8#0657# => '0' & O"054",
    8#0660# => '1' & O"247",
    8#0661# => '0' & O"267",
    8#0662# => '0' & O"742",
    8#0663# => '1' & O"426",
    8#0664# => '1' & O"313",
    8#0665# => '1' & O"626",
    8#0666# => '0' & O"426",
    8#0667# => '0' & O"034",
    8#0670# => '0' & O"054",
    8#0671# => '1' & O"317",
    8#0672# => '0' & O"267",
    8#0673# => '0' & O"034",
    8#0674# => '1' & O"626",
    8#0675# => '1' & O"557",
    8#0676# => '0' & O"020",
    8#0677# => '0' & O"572",
    8#0700# => '0' & O"572",
    8#0701# => '1' & O"352",
    8#0702# => '1' & O"536",
    8#0703# => '1' & O"176",
    8#0704# => '1' & O"433",
    8#0705# => '0' & O"420",
    8#0706# => '1' & O"006",
    8#0707# => '1' & O"453",
    8#0710# => '0' & O"376",
    8#0711# => '1' & O"456",
    8#0712# => '1' & O"416",
    8#0713# => '0' & O"420",
    8#0714# => '0' & O"316",
    8#0715# => '1' & O"314",
    8#0716# => '0' & O"730",
    8#0717# => '1' & O"030",
    8#0720# => '0' & O"530",
    8#0721# => '0' & O"330",
    8#0722# => '1' & O"130",
    8#0723# => '1' & O"030",
    8#0724# => '0' & O"130",
    8#0725# => '0' & O"630",
    8#0726# => '0' & O"330",
    8#0727# => '0' & O"530",
    8#0730# => '1' & O"414",
    8#0731# => '0' & O"060",
    8#0732# => '0' & O"020",
    8#0733# => '1' & O"612",
    8#0734# => '1' & O"573",
    8#0735# => '0' & O"542",
    8#0736# => '0' & O"776",
    8#0737# => '0' & O"054",
    8#0740# => '1' & O"357",
    8#0741# => '1' & O"652",
    8#0742# => '1' & O"352",
    8#0743# => '0' & O"142",
    8#0744# => '1' & O"633",
    8#0745# => '1' & O"316",
    8#0746# => '1' & O"116",
    8#0747# => '1' & O"052",
    8#0750# => '0' & O"312",
    8#0751# => '1' & O"414",
    8#0752# => '1' & O"273",
    8#0753# => '0' & O"420",
    8#0754# => '1' & O"222",
    8#0755# => '1' & O"222",
    8#0756# => '0' & O"576",
    8#0757# => '1' & O"663",
    8#0760# => '0' & O"722",
    8#0761# => '1' & O"422",
    8#0762# => '1' & O"062",
    8#0763# => '0' & O"216",
    8#0764# => '1' & O"576",
    8#0765# => '1' & O"673",
    8#0766# => '1' & O"662",
    8#0767# => '0' & O"650",
    8#0770# => '0' & O"036",
    8#0771# => '0' & O"007",
    8#0772# => '0' & O"416",
    8#0773# => '1' & O"662",
    8#0774# => '0' & O"450",
    8#0775# => '1' & O"222",
    8#0776# => '0' & O"576",
    8#0777# => '1' & O"076",
    8#1000# => '0' & O"020",
    8#1001# => '1' & O"476",
    8#1002# => '1' & O"776",
    8#1003# => '1' & O"126",
    8#1004# => '0' & O"422",
    8#1005# => '0' & O"113",
    8#1006# => '0' & O"650",
    8#1007# => '1' & O"231",
    8#1010# => '0' & O"616",
    8#1011# => '1' & O"024",
    8#1012# => '0' & O"413",
    8#1013# => '1' & O"356",
    8#1014# => '1' & O"506",
    8#1015# => '0' & O"003",
    8#1016# => '1' & O"316",
    8#1017# => '0' & O"576",
    8#1020# => '0' & O"003",
    8#1021# => '0' & O"776",
    8#1022# => '0' & O"456",
    8#1023# => '1' & O"131",
    8#1024# => '1' & O"542",
    8#1025# => '0' & O"107",
    8#1026# => '1' & O"462",
    8#1027# => '1' & O"636",
    8#1030# => '0' & O"007",
    8#1031# => '0' & O"714",
    8#1032# => '0' & O"665",
    8#1033# => '1' & O"014",
    8#1034# => '1' & O"165",
    8#1035# => '1' & O"114",
    8#1036# => '1' & O"161",
    8#1037# => '1' & O"771",
    8#1040# => '1' & O"214",
    8#1041# => '1' & O"161",
    8#1042# => '0' & O"765",
    8#1043# => '1' & O"314",
    8#1044# => '1' & O"161",
    8#1045# => '1' & O"575",
    8#1046# => '1' & O"161",
    8#1047# => '1' & O"345",
    8#1050# => '1' & O"161",
    8#1051# => '1' & O"731",
    8#1052# => '1' & O"656",
    8#1053# => '0' & O"516",
    8#1054# => '0' & O"032",
    8#1055# => '0' & O"277",
    8#1056# => '0' & O"516",
    8#1057# => '1' & O"456",
    8#1060# => '0' & O"034",
    8#1061# => '0' & O"416",
    8#1062# => '0' & O"154",
    8#1063# => '0' & O"303",
    8#1064# => '1' & O"656",
    8#1065# => '0' & O"676",
    8#1066# => '0' & O"343",
    8#1067# => '0' & O"346",
    8#1070# => '0' & O"752",
    8#1071# => '1' & O"314",
    8#1072# => '1' & O"425",
    8#1073# => '1' & O"124",
    8#1074# => '0' & O"033",
    8#1075# => '0' & O"524",
    8#1076# => '1' & O"123",
    8#1077# => '1' & O"731",
    8#1100# => '1' & O"235",
    8#1101# => '1' & O"123",
    8#1102# => '1' & O"731",
    8#1103# => '1' & O"661",
    8#1104# => '1' & O"345",
    8#1105# => '1' & O"314",
    8#1106# => '1' & O"155",
    8#1107# => '1' & O"575",
    8#1110# => '1' & O"214",
    8#1111# => '1' & O"155",
    8#1112# => '0' & O"765",
    8#1113# => '1' & O"114",
    8#1114# => '1' & O"155",
    8#1115# => '1' & O"771",
    8#1116# => '1' & O"014",
    8#1117# => '1' & O"155",
    8#1120# => '1' & O"155",
    8#1121# => '1' & O"155",
    8#1122# => '0' & O"614",
    8#1123# => '1' & O"362",
    8#1124# => '1' & O"514",
    8#1125# => '1' & O"056",
    8#1126# => '1' & O"656",
    8#1127# => '0' & O"630",
    8#1130# => '1' & O"073",
    8#1131# => '0' & O"224",
    8#1132# => '0' & O"573",
    8#1133# => '1' & O"752",
    8#1134# => '1' & O"172",
    8#1135# => '1' & O"413",
    8#1136# => '1' & O"426",
    8#1137# => '0' & O"547",
    8#1140# => '1' & O"626",
    8#1141# => '0' & O"416",
    8#1142# => '0' & O"552",
    8#1143# => '0' & O"563",
    8#1144# => '1' & O"316",
    8#1145# => '0' & O"322",
    8#1146# => '1' & O"652",
    8#1147# => '0' & O"676",
    8#1150# => '0' & O"663",
    8#1151# => '1' & O"456",
    8#1152# => '1' & O"416",
    8#1153# => '0' & O"356",
    8#1154# => '1' & O"316",
    8#1155# => '1' & O"056",
    8#1156# => '0' & O"316",
    8#1157# => '0' & O"546",
    8#1160# => '0' & O"224",
    8#1161# => '0' & O"733",
    8#1162# => '0' & O"430",
    8#1163# => '0' & O"746",
    8#1164# => '0' & O"747",
    8#1165# => '0' & O"630",
    8#1166# => '0' & O"154",
    8#1167# => '0' & O"727",
    8#1170# => '1' & O"116",
    8#1171# => '1' & O"116",
    8#1172# => '0' & O"224",
    8#1173# => '1' & O"123",
    8#1174# => '0' & O"060",
    8#1175# => '0' & O"714",
    8#1176# => '0' & O"330",
    8#1177# => '0' & O"330",
    8#1200# => '0' & O"030",
    8#1201# => '1' & O"030",
    8#1202# => '0' & O"530",
    8#1203# => '0' & O"030",
    8#1204# => '1' & O"130",
    8#1205# => '1' & O"653",
    8#1206# => '1' & O"131",
    8#1207# => '1' & O"742",
    8#1210# => '0' & O"456",
    8#1211# => '0' & O"576",
    8#1212# => '1' & O"033",
    8#1213# => '1' & O"322",
    8#1214# => '1' & O"656",
    8#1215# => '0' & O"426",
    8#1216# => '1' & O"656",
    8#1217# => '1' & O"576",
    8#1220# => '1' & O"043",
    8#1221# => '1' & O"456",
    8#1222# => '1' & O"742",
    8#1223# => '1' & O"461",
    8#1224# => '0' & O"220",
    8#1225# => '1' & O"322",
    8#1226# => '1' & O"576",
    8#1227# => '1' & O"127",
    8#1230# => '1' & O"376",
    8#1231# => '1' & O"616",
    8#1232# => '0' & O"060",
    8#1233# => '0' & O"220",
    8#1234# => '1' & O"316",
    8#1235# => '1' & O"056",
    8#1236# => '1' & O"203",
    8#1237# => '1' & O"616",
    8#1240# => '0' & O"576",
    8#1241# => '1' & O"177",
    8#1242# => '1' & O"656",
    8#1243# => '0' & O"426",
    8#1244# => '1' & O"656",
    8#1245# => '0' & O"667",
    8#1246# => '0' & O"314",
    8#1247# => '0' & O"712",
    8#1250# => '0' & O"536",
    8#1251# => '1' & O"257",
    8#1252# => '0' & O"276",
    8#1253# => '1' & O"446",
    8#1254# => '1' & O"356",
    8#1255# => '1' & O"454",
    8#1256# => '1' & O"427",
    8#1257# => '0' & O"146",
    8#1260# => '1' & O"333",
    8#1261# => '0' & O"124",
    8#1262# => '0' & O"003",
    8#1263# => '0' & O"222",
    8#1264# => '1' & O"546",
    8#1265# => '0' & O"772",
    8#1266# => '1' & O"062",
    8#1267# => '1' & O"646",
    8#1270# => '0' & O"220",
    8#1271# => '1' & O"044",
    8#1272# => '0' & O"630",
    8#1273# => '1' & O"130",
    8#1274# => '0' & O"330",
    8#1275# => '0' & O"130",
    8#1276# => '0' & O"430",
    8#1277# => '0' & O"730",
    8#1300# => '0' & O"130",
    8#1301# => '1' & O"633",
    8#1302# => '1' & O"746",
    8#1303# => '0' & O"623",
    8#1304# => '1' & O"616",
    8#1305# => '0' & O"542",
    8#1306# => '1' & O"423",
    8#1307# => '1' & O"316",
    8#1310# => '0' & O"074",
    8#1311# => '1' & O"554",
    8#1312# => '1' & O"427",
    8#1313# => '0' & O"752",
    8#1314# => '1' & O"376",
    8#1315# => '1' & O"414",
    8#1316# => '0' & O"056",
    8#1317# => '1' & O"142",
    8#1320# => '1' & O"533",
    8#1321# => '0' & O"416",
    8#1322# => '0' & O"552",
    8#1323# => '1' & O"156",
    8#1324# => '1' & O"477",
    8#1325# => '0' & O"316",
    8#1326# => '0' & O"452",
    8#1327# => '1' & O"616",
    8#1330# => '1' & O"176",
    8#1331# => '1' & O"437",
    8#1332# => '1' & O"646",
    8#1333# => '0' & O"616",
    8#1334# => '0' & O"056",
    8#1335# => '1' & O"414",
    8#1336# => '0' & O"753",
    8#1337# => '1' & O"114",
    8#1340# => '0' & O"330",
    8#1341# => '0' & O"130",
    8#1342# => '0' & O"030",
    8#1343# => '0' & O"130",
    8#1344# => '0' & O"730",
    8#1345# => '1' & O"130",
    8#1346# => '1' & O"030",
    8#1347# => '0' & O"030",
    8#1350# => '0' & O"530",
    8#1351# => '0' & O"530",
    8#1352# => '0' & O"330",
    8#1353# => '1' & O"567",
    8#1354# => '1' & O"656",
    8#1355# => '0' & O"456",
    8#1356# => '0' & O"606",
    8#1357# => '1' & O"272",
    8#1360# => '0' & O"573",
    8#1361# => '0' & O"772",
    8#1362# => '1' & O"316",
    8#1363# => '0' & O"752",
    8#1364# => '1' & O"713",
    8#1365# => '0' & O"637",
    8#1366# => '0' & O"316",
    8#1367# => '1' & O"414",
    8#1370# => '0' & O"230",
    8#1371# => '0' & O"330",
    8#1372# => '0' & O"030",
    8#1373# => '0' & O"230",
    8#1374# => '0' & O"530",
    8#1375# => '1' & O"007",
    8#1376# => '0' & O"514",
    8#1377# => '0' & O"773"
  );

  constant ROM_45 : RomType := (
    8#0000# => '0' & O"255",
    8#0001# => '1' & O"420",
    8#0002# => '0' & O"451",
    8#0003# => '1' & O"456",
    8#0004# => '1' & O"746",
    8#0005# => '0' & O"472",
    8#0006# => '1' & O"572",
    8#0007# => '1' & O"616",
    8#0010# => '1' & O"352",
    8#0011# => '1' & O"611",
    8#0012# => '1' & O"611",
    8#0013# => '1' & O"352",
    8#0014# => '1' & O"445",
    8#0015# => '0' & O"623",
    8#0016# => '1' & O"024",
    8#0017# => '0' & O"507",
    8#0020# => '1' & O"035",
    8#0021# => '1' & O"656",
    8#0022# => '0' & O"616",
    8#0023# => '0' & O"013",
    8#0024# => '1' & O"220",
    8#0025# => '1' & O"035",
    8#0026# => '1' & O"656",
    8#0027# => '1' & O"020",
    8#0030# => '0' & O"220",
    8#0031# => '0' & O"324",
    8#0032# => '0' & O"143",
    8#0033# => '0' & O"450",
    8#0034# => '0' & O"316",
    8#0035# => '1' & O"160",
    8#0036# => '0' & O"000",
    8#0037# => '1' & O"370",
    8#0040# => '1' & O"656",
    8#0041# => '1' & O"171",
    8#0042# => '1' & O"431",
    8#0043# => '1' & O"211",
    8#0044# => '1' & O"431",
    8#0045# => '1' & O"376",
    8#0046# => '1' & O"370",
    8#0047# => '0' & O"676",
    8#0050# => '0' & O"267",
    8#0051# => '1' & O"576",
    8#0052# => '0' & O"265",
    8#0053# => '0' & O"123",
    8#0054# => '0' & O"220",
    8#0055# => '1' & O"656",
    8#0056# => '1' & O"024",
    8#0057# => '1' & O"713",
    8#0060# => '0' & O"376",
    8#0061# => '1' & O"711",
    8#0062# => '0' & O"124",
    8#0063# => '0' & O"263",
    8#0064# => '1' & O"224",
    8#0065# => '0' & O"647",
    8#0066# => '0' & O"353",
    8#0067# => '0' & O"220",
    8#0070# => '0' & O"616",
    8#0071# => '0' & O"220",
    8#0072# => '1' & O"656",
    8#0073# => '0' & O"616",
    8#0074# => '0' & O"772",
    8#0075# => '0' & O"433",
    8#0076# => '0' & O"652",
    8#0077# => '0' & O"433",
    8#0100# => '0' & O"316",
    8#0101# => '0' & O"014",
    8#0102# => '0' & O"530",
    8#0103# => '1' & O"414",
    8#0104# => '0' & O"712",
    8#0105# => '1' & O"657",
    8#0106# => '1' & O"224",
    8#0107# => '0' & O"727",
    8#0110# => '1' & O"656",
    8#0111# => '0' & O"343",
    8#0112# => '0' & O"312",
    8#0113# => '0' & O"014",
    8#0114# => '0' & O"530",
    8#0115# => '1' & O"512",
    8#0116# => '1' & O"172",
    8#0117# => '1' & O"463",
    8#0120# => '1' & O"777",
    8#0121# => '0' & O"451",
    8#0122# => '1' & O"615",
    8#0123# => '0' & O"056",
    8#0124# => '1' & O"462",
    8#0125# => '1' & O"456",
    8#0126# => '0' & O"416",
    8#0127# => '1' & O"625",
    8#0130# => '0' & O"704",
    8#0131# => '1' & O"445",
    8#0132# => '0' & O"316",
    8#0133# => '0' & O"330",
    8#0134# => '0' & O"630",
    8#0135# => '1' & O"414",
    8#0136# => '1' & O"171",
    8#0137# => '1' & O"031",
    8#0140# => '0' & O"767",
    8#0141# => '0' & O"752",
    8#0142# => '0' & O"742",
    8#0143# => '1' & O"017",
    8#0144# => '0' & O"316",
    8#0145# => '0' & O"214",
    8#0146# => '0' & O"430",
    8#0147# => '1' & O"656",
    8#0150# => '0' & O"007",
    8#0151# => '0' & O"220",
    8#0152# => '0' & O"704",
    8#0153# => '0' & O"424",
    8#0154# => '0' & O"717",
    8#0155# => '1' & O"256",
    8#0156# => '0' & O"736",
    8#0157# => '1' & O"146",
    8#0160# => '0' & O"713",
    8#0161# => '0' & O"376",
    8#0162# => '1' & O"231",
    8#0163# => '0' & O"104",
    8#0164# => '0' & O"127",
    8#0165# => '0' & O"220",
    8#0166# => '1' & O"024",
    8#0167# => '0' & O"653",
    8#0170# => '1' & O"035",
    8#0171# => '0' & O"104",
    8#0172# => '1' & O"224",
    8#0173# => '0' & O"353",
    8#0174# => '1' & O"717",
    8#0175# => '1' & O"656",
    8#0176# => '0' & O"620",
    8#0177# => '0' & O"552",
    8#0200# => '0' & O"552",
    8#0201# => '0' & O"704",
    8#0202# => '0' & O"542",
    8#0203# => '1' & O"224",
    8#0204# => '1' & O"173",
    8#0205# => '1' & O"213",
    8#0206# => '1' & O"244",
    8#0207# => '0' & O"704",
    8#0210# => '0' & O"444",
    8#0211# => '0' & O"604",
    8#0212# => '1' & O"250",
    8#0213# => '0' & O"676",
    8#0214# => '1' & O"073",
    8#0215# => '0' & O"404",
    8#0216# => '0' & O"776",
    8#0217# => '1' & O"107",
    8#0220# => '0' & O"644",
    8#0221# => '0' & O"316",
    8#0222# => '0' & O"752",
    8#0223# => '0' & O"124",
    8#0224# => '1' & O"403",
    8#0225# => '0' & O"424",
    8#0226# => '1' & O"607",
    8#0227# => '0' & O"744",
    8#0230# => '0' & O"624",
    8#0231# => '1' & O"013",
    8#0232# => '0' & O"607",
    8#0233# => '1' & O"253",
    8#0234# => '1' & O"224",
    8#0235# => '1' & O"213",
    8#0236# => '1' & O"304",
    8#0237# => '0' & O"144",
    8#0240# => '0' & O"056",
    8#0241# => '1' & O"227",
    8#0242# => '1' & O"304",
    8#0243# => '0' & O"144",
    8#0244# => '0' & O"220",
    8#0245# => '0' & O"220",
    8#0246# => '1' & O"304",
    8#0247# => '0' & O"376",
    8#0250# => '0' & O"144",
    8#0251# => '0' & O"244",
    8#0252# => '0' & O"056",
    8#0253# => '1' & O"772",
    8#0254# => '1' & O"772",
    8#0255# => '0' & O"772",
    8#0256# => '0' & O"772",
    8#0257# => '0' & O"112",
    8#0260# => '1' & O"313",
    8#0261# => '1' & O"656",
    8#0262# => '1' & O"646",
    8#0263# => '0' & O"646",
    8#0264# => '1' & O"333",
    8#0265# => '1' & O"656",
    8#0266# => '1' & O"046",
    8#0267# => '0' & O"112",
    8#0270# => '1' & O"373",
    8#0271# => '1' & O"216",
    8#0272# => '1' & O"752",
    8#0273# => '0' & O"016",
    8#0274# => '1' & O"373",
    8#0275# => '1' & O"337",
    8#0276# => '0' & O"220",
    8#0277# => '1' & O"777",
    8#0300# => '0' & O"624",
    8#0301# => '1' & O"607",
    8#0302# => '0' & O"744",
    8#0303# => '0' & O"424",
    8#0304# => '1' & O"013",
    8#0305# => '0' & O"777",
    8#0306# => '0' & O"650",
    8#0307# => '0' & O"450",
    8#0310# => '0' & O"060",
    8#0311# => '1' & O"304",
    8#0312# => '0' & O"220",
    8#0313# => '0' & O"220",
    8#0314# => '1' & O"046",
    8#0315# => '1' & O"216",
    8#0316# => '1' & O"752",
    8#0317# => '1' & O"467",
    8#0320# => '1' & O"356",
    8#0321# => '0' & O"614",
    8#0322# => '0' & O"060",
    8#0323# => '1' & O"324",
    8#0324# => '1' & O"543",
    8#0325# => '1' & O"256",
    8#0326# => '0' & O"704",
    8#0327# => '1' & O"163",
    8#0330# => '0' & O"220",
    8#0331# => '1' & O"414",
    8#0332# => '1' & O"517",
    8#0333# => '1' & O"324",
    8#0334# => '1' & O"747",
    8#0335# => '1' & O"304",
    8#0336# => '0' & O"724",
    8#0337# => '1' & O"457",
    8#0340# => '1' & O"344",
    8#0341# => '0' & O"060",
    8#0342# => '0' & O"056",
    8#0343# => '1' & O"462",
    8#0344# => '1' & O"216",
    8#0345# => '1' & O"214",
    8#0346# => '1' & O"616",
    8#0347# => '0' & O"034",
    8#0350# => '0' & O"454",
    8#0351# => '1' & O"633",
    8#0352# => '0' & O"060",
    8#0353# => '0' & O"316",
    8#0354# => '0' & O"742",
    8#0355# => '1' & O"224",
    8#0356# => '0' & O"337",
    8#0357# => '0' & O"647",
    8#0360# => '0' & O"124",
    8#0361# => '0' & O"773",
    8#0362# => '1' & O"656",
    8#0363# => '0' & O"316",
    8#0364# => '0' & O"542",
    8#0365# => '1' & O"160",
    8#0366# => '0' & O"316",
    8#0367# => '1' & O"360",
    8#0370# => '0' & O"767",
    8#0371# => '0' & O"324",
    8#0372# => '1' & O"703",
    8#0373# => '1' & O"224",
    8#0374# => '1' & O"773",
    8#0375# => '1' & O"020",
    8#0376# => '1' & O"220",
    8#0377# => '0' & O"420",
    8#0400# => '1' & O"076",
    8#0401# => '1' & O"717",
    8#0402# => '1' & O"456",
    8#0403# => '0' & O"301",
    8#0404# => '1' & O"370",
    8#0405# => '1' & O"656",
    8#0406# => '0' & O"301",
    8#0407# => '1' & O"370",
    8#0410# => '1' & O"656",
    8#0411# => '1' & O"124",
    8#0412# => '0' & O"063",
    8#0413# => '1' & O"656",
    8#0414# => '0' & O"524",
    8#0415# => '0' & O"153",
    8#0416# => '0' & O"176",
    8#0417# => '0' & O"107",
    8#0420# => '1' & O"044",
    8#0421# => '0' & O"336",
    8#0422# => '1' & O"231",
    8#0423# => '1' & O"360",
    8#0424# => '1' & O"225",
    8#0425# => '1' & O"141",
    8#0426# => '0' & O"265",
    8#0427# => '1' & O"370",
    8#0430# => '0' & O"020",
    8#0431# => '1' & O"656",
    8#0432# => '1' & O"231",
    8#0433# => '1' & O"224",
    8#0434# => '1' & O"553",
    8#0435# => '1' & O"356",
    8#0436# => '1' & O"742",
    8#0437# => '0' & O"446",
    8#0440# => '1' & O"646",
    8#0441# => '0' & O"552",
    8#0442# => '1' & O"222",
    8#0443# => '0' & O"672",
    8#0444# => '0' & O"207",
    8#0445# => '1' & O"322",
    8#0446# => '0' & O"752",
    8#0447# => '0' & O"227",
    8#0450# => '1' & O"316",
    8#0451# => '1' & O"216",
    8#0452# => '1' & O"360",
    8#0453# => '1' & O"056",
    8#0454# => '0' & O"433",
    8#0455# => '1' & O"056",
    8#0456# => '0' & O"414",
    8#0457# => '1' & O"573",
    8#0460# => '1' & O"360",
    8#0461# => '1' & O"656",
    8#0462# => '0' & O"642",
    8#0463# => '0' & O"327",
    8#0464# => '0' & O"256",
    8#0465# => '0' & O"616",
    8#0466# => '0' & O"212",
    8#0467# => '1' & O"457",
    8#0470# => '0' & O"047",
    8#0471# => '0' & O"020",
    8#0472# => '0' & O"524",
    8#0473# => '0' & O"167",
    8#0474# => '0' & O"376",
    8#0475# => '1' & O"676",
    8#0476# => '0' & O"117",
    8#0477# => '1' & O"222",
    8#0500# => '1' & O"576",
    8#0501# => '0' & O"377",
    8#0502# => '0' & O"776",
    8#0503# => '1' & O"462",
    8#0504# => '0' & O"722",
    8#0505# => '1' & O"456",
    8#0506# => '0' & O"456",
    8#0507# => '1' & O"522",
    8#0510# => '0' & O"403",
    8#0511# => '1' & O"656",
    8#0512# => '1' & O"370",
    8#0513# => '1' & O"116",
    8#0514# => '1' & O"676",
    8#0515# => '1' & O"456",
    8#0516# => '0' & O"422",
    8#0517# => '1' & O"360",
    8#0520# => '1' & O"776",
    8#0521# => '1' & O"776",
    8#0522# => '0' & O"257",
    8#0523# => '0' & O"316",
    8#0524# => '0' & O"052",
    8#0525# => '1' & O"326",
    8#0526# => '1' & O"311",
    8#0527# => '1' & O"542",
    8#0530# => '1' & O"370",
    8#0531# => '0' & O"414",
    8#0532# => '1' & O"221",
    8#0533# => '0' & O"614",
    8#0534# => '1' & O"155",
    8#0535# => '1' & O"014",
    8#0536# => '1' & O"155",
    8#0537# => '0' & O"214",
    8#0540# => '1' & O"030",
    8#0541# => '1' & O"214",
    8#0542# => '1' & O"155",
    8#0543# => '1' & O"071",
    8#0544# => '1' & O"155",
    8#0545# => '1' & O"461",
    8#0546# => '0' & O"416",
    8#0547# => '1' & O"155",
    8#0550# => '0' & O"216",
    8#0551# => '1' & O"455",
    8#0552# => '1' & O"461",
    8#0553# => '1' & O"256",
    8#0554# => '1' & O"224",
    8#0555# => '0' & O"727",
    8#0556# => '1' & O"124",
    8#0557# => '0' & O"727",
    8#0560# => '1' & O"656",
    8#0561# => '0' & O"376",
    8#0562# => '1' & O"151",
    8#0563# => '1' & O"461",
    8#0564# => '1' & O"256",
    8#0565# => '0' & O"020",
    8#0566# => '1' & O"461",
    8#0567# => '1' & O"256",
    8#0570# => '1' & O"256",
    8#0571# => '1' & O"125",
    8#0572# => '1' & O"256",
    8#0573# => '1' & O"655",
    8#0574# => '1' & O"461",
    8#0575# => '1' & O"214",
    8#0576# => '1' & O"161",
    8#0577# => '1' & O"071",
    8#0600# => '1' & O"014",
    8#0601# => '1' & O"165",
    8#0602# => '0' & O"214",
    8#0603# => '1' & O"030",
    8#0604# => '0' & O"614",
    8#0605# => '1' & O"161",
    8#0606# => '0' & O"414",
    8#0607# => '1' & O"161",
    8#0610# => '1' & O"161",
    8#0611# => '1' & O"456",
    8#0612# => '1' & O"116",
    8#0613# => '1' & O"514",
    8#0614# => '0' & O"530",
    8#0615# => '1' & O"763",
    8#0616# => '0' & O"614",
    8#0617# => '1' & O"030",
    8#0620# => '0' & O"630",
    8#0621# => '0' & O"530",
    8#0622# => '0' & O"230",
    8#0623# => '0' & O"430",
    8#0624# => '1' & O"130",
    8#0625# => '0' & O"124",
    8#0626# => '1' & O"553",
    8#0627# => '0' & O"060",
    8#0630# => '1' & O"356",
    8#0631# => '1' & O"742",
    8#0632# => '0' & O"020",
    8#0633# => '0' & O"420",
    8#0634# => '0' & O"416",
    8#0635# => '1' & O"226",
    8#0636# => '1' & O"056",
    8#0637# => '1' & O"207",
    8#0640# => '0' & O"776",
    8#0641# => '1' & O"416",
    8#0642# => '1' & O"203",
    8#0643# => '1' & O"616",
    8#0644# => '0' & O"420",
    8#0645# => '0' & O"420",
    8#0646# => '0' & O"512",
    8#0647# => '0' & O"420",
    8#0650# => '0' & O"742",
    8#0651# => '1' & O"516",
    8#0652# => '1' & O"243",
    8#0653# => '1' & O"716",
    8#0654# => '0' & O"416",
    8#0655# => '0' & O"034",
    8#0656# => '1' & O"122",
    8#0657# => '0' & O"054",
    8#0660# => '1' & O"247",
    8#0661# => '0' & O"327",
    8#0662# => '0' & O"742",
    8#0663# => '1' & O"426",
    8#0664# => '1' & O"313",
    8#0665# => '1' & O"626",
    8#0666# => '0' & O"426",
    8#0667# => '0' & O"034",
    8#0670# => '0' & O"054",
    8#0671# => '1' & O"317",
    8#0672# => '0' & O"327",
    8#0673# => '0' & O"034",
    8#0674# => '1' & O"626",
    8#0675# => '1' & O"557",
    8#0676# => '0' & O"020",
    8#0677# => '0' & O"572",
    8#0700# => '0' & O"572",
    8#0701# => '1' & O"352",
    8#0702# => '1' & O"536",
    8#0703# => '1' & O"176",
    8#0704# => '1' & O"433",
    8#0705# => '0' & O"420",
    8#0706# => '1' & O"006",
    8#0707# => '1' & O"453",
    8#0710# => '0' & O"376",
    8#0711# => '1' & O"456",
    8#0712# => '1' & O"416",
    8#0713# => '0' & O"420",
    8#0714# => '0' & O"316",
    8#0715# => '1' & O"314",
    8#0716# => '0' & O"730",
    8#0717# => '1' & O"030",
    8#0720# => '0' & O"530",
    8#0721# => '0' & O"330",
    8#0722# => '1' & O"130",
    8#0723# => '1' & O"030",
    8#0724# => '0' & O"130",
    8#0725# => '0' & O"630",
    8#0726# => '0' & O"330",
    8#0727# => '0' & O"530",
    8#0730# => '0' & O"020",
    8#0731# => '0' & O"060",
    8#0732# => '0' & O"020",
    8#0733# => '1' & O"612",
    8#0734# => '1' & O"573",
    8#0735# => '0' & O"542",
    8#0736# => '0' & O"776",
    8#0737# => '0' & O"054",
    8#0740# => '1' & O"357",
    8#0741# => '1' & O"652",
    8#0742# => '1' & O"352",
    8#0743# => '0' & O"142",
    8#0744# => '1' & O"633",
    8#0745# => '1' & O"316",
    8#0746# => '1' & O"116",
    8#0747# => '1' & O"052",
    8#0750# => '0' & O"312",
    8#0751# => '1' & O"414",
    8#0752# => '1' & O"273",
    8#0753# => '0' & O"420",
    8#0754# => '1' & O"222",
    8#0755# => '1' & O"222",
    8#0756# => '0' & O"576",
    8#0757# => '1' & O"663",
    8#0760# => '0' & O"722",
    8#0761# => '1' & O"422",
    8#0762# => '1' & O"062",
    8#0763# => '0' & O"216",
    8#0764# => '1' & O"576",
    8#0765# => '1' & O"673",
    8#0766# => '1' & O"676",
    8#0767# => '1' & O"370",
    8#0770# => '1' & O"656",
    8#0771# => '0' & O"036",
    8#0772# => '0' & O"013",
    8#0773# => '0' & O"416",
    8#0774# => '1' & O"662",
    8#0775# => '1' & O"360",
    8#0776# => '1' & O"222",
    8#0777# => '0' & O"576",
    8#1000# => '1' & O"420",
    8#1001# => '1' & O"476",
    8#1002# => '1' & O"776",
    8#1003# => '1' & O"126",
    8#1004# => '0' & O"422",
    8#1005# => '0' & O"113",
    8#1006# => '0' & O"650",
    8#1007# => '1' & O"231",
    8#1010# => '0' & O"616",
    8#1011# => '1' & O"024",
    8#1012# => '0' & O"413",
    8#1013# => '1' & O"356",
    8#1014# => '1' & O"506",
    8#1015# => '0' & O"003",
    8#1016# => '1' & O"316",
    8#1017# => '0' & O"576",
    8#1020# => '0' & O"003",
    8#1021# => '0' & O"776",
    8#1022# => '0' & O"456",
    8#1023# => '1' & O"131",
    8#1024# => '1' & O"542",
    8#1025# => '0' & O"107",
    8#1026# => '1' & O"462",
    8#1027# => '1' & O"636",
    8#1030# => '0' & O"007",
    8#1031# => '0' & O"714",
    8#1032# => '0' & O"665",
    8#1033# => '1' & O"014",
    8#1034# => '1' & O"165",
    8#1035# => '1' & O"114",
    8#1036# => '1' & O"161",
    8#1037# => '1' & O"771",
    8#1040# => '1' & O"214",
    8#1041# => '1' & O"161",
    8#1042# => '0' & O"765",
    8#1043# => '1' & O"314",
    8#1044# => '1' & O"161",
    8#1045# => '1' & O"575",
    8#1046# => '1' & O"161",
    8#1047# => '1' & O"345",
    8#1050# => '1' & O"161",
    8#1051# => '1' & O"731",
    8#1052# => '1' & O"656",
    8#1053# => '0' & O"516",
    8#1054# => '0' & O"032",
    8#1055# => '0' & O"277",
    8#1056# => '0' & O"516",
    8#1057# => '1' & O"456",
    8#1060# => '0' & O"034",
    8#1061# => '0' & O"416",
    8#1062# => '0' & O"154",
    8#1063# => '0' & O"303",
    8#1064# => '1' & O"656",
    8#1065# => '0' & O"676",
    8#1066# => '0' & O"343",
    8#1067# => '0' & O"346",
    8#1070# => '0' & O"752",
    8#1071# => '1' & O"314",
    8#1072# => '1' & O"425",
    8#1073# => '1' & O"124",
    8#1074# => '0' & O"033",
    8#1075# => '0' & O"524",
    8#1076# => '1' & O"123",
    8#1077# => '1' & O"731",
    8#1100# => '1' & O"235",
    8#1101# => '1' & O"123",
    8#1102# => '1' & O"731",
    8#1103# => '1' & O"661",
    8#1104# => '1' & O"345",
    8#1105# => '1' & O"314",
    8#1106# => '1' & O"155",
    8#1107# => '1' & O"575",
    8#1110# => '1' & O"214",
    8#1111# => '1' & O"155",
    8#1112# => '0' & O"765",
    8#1113# => '1' & O"114",
    8#1114# => '1' & O"155",
    8#1115# => '1' & O"771",
    8#1116# => '1' & O"014",
    8#1117# => '1' & O"155",
    8#1120# => '1' & O"155",
    8#1121# => '1' & O"155",
    8#1122# => '0' & O"614",
    8#1123# => '1' & O"362",
    8#1124# => '1' & O"514",
    8#1125# => '1' & O"056",
    8#1126# => '1' & O"656",
    8#1127# => '0' & O"630",
    8#1130# => '1' & O"073",
    8#1131# => '0' & O"224",
    8#1132# => '0' & O"573",
    8#1133# => '1' & O"752",
    8#1134# => '1' & O"172",
    8#1135# => '1' & O"413",
    8#1136# => '1' & O"426",
    8#1137# => '0' & O"547",
    8#1140# => '1' & O"626",
    8#1141# => '0' & O"416",
    8#1142# => '0' & O"552",
    8#1143# => '0' & O"563",
    8#1144# => '1' & O"316",
    8#1145# => '0' & O"322",
    8#1146# => '1' & O"652",
    8#1147# => '0' & O"676",
    8#1150# => '0' & O"663",
    8#1151# => '1' & O"456",
    8#1152# => '1' & O"416",
    8#1153# => '0' & O"356",
    8#1154# => '1' & O"316",
    8#1155# => '1' & O"056",
    8#1156# => '0' & O"316",
    8#1157# => '0' & O"546",
    8#1160# => '0' & O"224",
    8#1161# => '0' & O"733",
    8#1162# => '0' & O"430",
    8#1163# => '0' & O"746",
    8#1164# => '0' & O"747",
    8#1165# => '0' & O"630",
    8#1166# => '0' & O"154",
    8#1167# => '0' & O"727",
    8#1170# => '1' & O"116",
    8#1171# => '1' & O"116",
    8#1172# => '0' & O"224",
    8#1173# => '1' & O"123",
    8#1174# => '0' & O"060",
    8#1175# => '0' & O"714",
    8#1176# => '0' & O"330",
    8#1177# => '0' & O"330",
    8#1200# => '0' & O"030",
    8#1201# => '1' & O"030",
    8#1202# => '0' & O"530",
    8#1203# => '0' & O"030",
    8#1204# => '1' & O"130",
    8#1205# => '1' & O"653",
    8#1206# => '1' & O"131",
    8#1207# => '1' & O"742",
    8#1210# => '0' & O"456",
    8#1211# => '0' & O"576",
    8#1212# => '1' & O"033",
    8#1213# => '1' & O"322",
    8#1214# => '1' & O"656",
    8#1215# => '0' & O"426",
    8#1216# => '1' & O"656",
    8#1217# => '1' & O"576",
    8#1220# => '1' & O"043",
    8#1221# => '1' & O"456",
    8#1222# => '1' & O"742",
    8#1223# => '1' & O"461",
    8#1224# => '0' & O"220",
    8#1225# => '1' & O"322",
    8#1226# => '1' & O"576",
    8#1227# => '1' & O"127",
    8#1230# => '1' & O"376",
    8#1231# => '1' & O"616",
    8#1232# => '0' & O"060",
    8#1233# => '0' & O"220",
    8#1234# => '1' & O"316",
    8#1235# => '1' & O"056",
    8#1236# => '1' & O"203",
    8#1237# => '1' & O"616",
    8#1240# => '0' & O"576",
    8#1241# => '1' & O"177",
    8#1242# => '1' & O"656",
    8#1243# => '0' & O"426",
    8#1244# => '1' & O"656",
    8#1245# => '0' & O"667",
    8#1246# => '0' & O"314",
    8#1247# => '0' & O"712",
    8#1250# => '0' & O"536",
    8#1251# => '1' & O"257",
    8#1252# => '0' & O"276",
    8#1253# => '1' & O"446",
    8#1254# => '1' & O"356",
    8#1255# => '1' & O"454",
    8#1256# => '1' & O"427",
    8#1257# => '0' & O"146",
    8#1260# => '1' & O"333",
    8#1261# => '0' & O"124",
    8#1262# => '0' & O"003",
    8#1263# => '1' & O"220",
    8#1264# => '1' & O"557",
    8#1265# => '0' & O"000",
    8#1266# => '1' & O"062",
    8#1267# => '1' & O"646",
    8#1270# => '0' & O"220",
    8#1271# => '1' & O"044",
    8#1272# => '0' & O"630",
    8#1273# => '1' & O"130",
    8#1274# => '0' & O"330",
    8#1275# => '0' & O"130",
    8#1276# => '0' & O"430",
    8#1277# => '0' & O"730",
    8#1300# => '0' & O"130",
    8#1301# => '1' & O"633",
    8#1302# => '1' & O"746",
    8#1303# => '0' & O"623",
    8#1304# => '1' & O"616",
    8#1305# => '0' & O"542",
    8#1306# => '1' & O"423",
    8#1307# => '1' & O"316",
    8#1310# => '0' & O"074",
    8#1311# => '1' & O"554",
    8#1312# => '1' & O"427",
    8#1313# => '0' & O"752",
    8#1314# => '1' & O"376",
    8#1315# => '1' & O"414",
    8#1316# => '0' & O"056",
    8#1317# => '1' & O"142",
    8#1320# => '1' & O"533",
    8#1321# => '0' & O"416",
    8#1322# => '0' & O"552",
    8#1323# => '1' & O"156",
    8#1324# => '1' & O"477",
    8#1325# => '0' & O"316",
    8#1326# => '0' & O"452",
    8#1327# => '1' & O"616",
    8#1330# => '1' & O"176",
    8#1331# => '1' & O"437",
    8#1332# => '1' & O"646",
    8#1333# => '0' & O"616",
    8#1334# => '0' & O"056",
    8#1335# => '1' & O"414",
    8#1336# => '0' & O"753",
    8#1337# => '1' & O"114",
    8#1340# => '0' & O"330",
    8#1341# => '0' & O"130",
    8#1342# => '0' & O"030",
    8#1343# => '0' & O"130",
    8#1344# => '0' & O"730",
    8#1345# => '1' & O"130",
    8#1346# => '1' & O"030",
    8#1347# => '0' & O"030",
    8#1350# => '0' & O"530",
    8#1351# => '0' & O"530",
    8#1352# => '0' & O"330",
    8#1353# => '1' & O"567",
    8#1354# => '1' & O"656",
    8#1355# => '0' & O"456",
    8#1356# => '0' & O"606",
    8#1357# => '1' & O"272",
    8#1360# => '0' & O"573",
    8#1361# => '0' & O"772",
    8#1362# => '1' & O"316",
    8#1363# => '0' & O"752",
    8#1364# => '1' & O"713",
    8#1365# => '0' & O"637",
    8#1366# => '0' & O"316",
    8#1367# => '1' & O"414",
    8#1370# => '0' & O"230",
    8#1371# => '0' & O"330",
    8#1372# => '0' & O"030",
    8#1373# => '0' & O"230",
    8#1374# => '0' & O"530",
    8#1375# => '1' & O"007",
    8#1376# => '0' & O"514",
    8#1377# => '0' & O"773",
    8#1400# => '1' & O"020",
    8#1401# => '0' & O"000",
    8#1402# => '0' & O"453",
    8#1403# => '0' & O"547",
    8#1404# => '0' & O"553",
    8#1405# => '0' & O"000",
    8#1406# => '0' & O"423",
    8#1407# => '0' & O"420",
    8#1410# => '1' & O"020",
    8#1411# => '1' & O"420",
    8#1412# => '0' & O"633",
    8#1413# => '0' & O"643",
    8#1414# => '1' & O"450",
    8#1415# => '0' & O"777",
    8#1416# => '0' & O"650",
    8#1417# => '0' & O"450",
    8#1420# => '0' & O"773",
    8#1421# => '0' & O"377",
    8#1422# => '1' & O"756",
    8#1423# => '1' & O"756",
    8#1424# => '1' & O"756",
    8#1425# => '0' & O"153",
    8#1426# => '1' & O"020",
    8#1427# => '1' & O"035",
    8#1430# => '0' & O"416",
    8#1431# => '0' & O"513",
    8#1432# => '1' & O"756",
    8#1433# => '1' & O"756",
    8#1434# => '1' & O"756",
    8#1435# => '0' & O"060",
    8#1436# => '1' & O"020",
    8#1437# => '0' & O"320",
    8#1440# => '1' & O"044",
    8#1441# => '1' & O"020",
    8#1442# => '0' & O"203",
    8#1443# => '0' & O"314",
    8#1444# => '0' & O"060",
    8#1445# => '1' & O"020",
    8#1446# => '0' & O"227",
    8#1447# => '0' & O"504",
    8#1450# => '0' & O"621",
    8#1451# => '0' & O"413",
    8#1452# => '0' & O"463",
    8#1453# => '0' & O"237",
    8#1454# => '1' & O"020",
    8#1455# => '0' & O"000",
    8#1456# => '0' & O"605",
    8#1457# => '0' & O"443",
    8#1460# => '0' & O"000",
    8#1461# => '0' & O"020",
    8#1462# => '1' & O"756",
    8#1463# => '1' & O"756",
    8#1464# => '1' & O"756",
    8#1465# => '0' & O"113",
    8#1466# => '1' & O"020",
    8#1467# => '0' & O"000",
    8#1470# => '1' & O"231",
    8#1471# => '1' & O"007",
    8#1472# => '1' & O"357",
    8#1473# => '1' & O"407",
    8#1474# => '0' & O"056",
    8#1475# => '1' & O"620",
    8#1476# => '0' & O"450",
    8#1477# => '1' & O"235",
    8#1500# => '1' & O"007",
    8#1501# => '0' & O"605",
    8#1502# => '1' & O"144",
    8#1503# => '0' & O"307",
    8#1504# => '0' & O"605",
    8#1505# => '1' & O"356",
    8#1506# => '1' & O"742",
    8#1507# => '0' & O"447",
    8#1510# => '1' & O"020",
    8#1511# => '1' & O"020",
    8#1512# => '1' & O"144",
    8#1513# => '0' & O"137",
    8#1514# => '0' & O"621",
    8#1515# => '1' & O"104",
    8#1516# => '0' & O"504",
    8#1517# => '0' & O"307",
    8#1520# => '0' & O"416",
    8#1521# => '1' & O"756",
    8#1522# => '0' & O"416",
    8#1523# => '0' & O"250",
    8#1524# => '1' & O"652",
    8#1525# => '0' & O"250",
    8#1526# => '0' & O"713",
    8#1527# => '0' & O"000",
    8#1530# => '0' & O"000",
    8#1531# => '1' & O"044",
    8#1532# => '1' & O"104",
    8#1533# => '0' & O"605",
    8#1534# => '0' & O"204",
    8#1535# => '0' & O"037",
    8#1536# => '1' & O"035",
    8#1537# => '0' & O"503",
    8#1540# => '0' & O"304",
    8#1541# => '1' & O"244",
    8#1542# => '1' & O"420",
    8#1543# => '1' & O"420",
    8#1544# => '0' & O"104",
    8#1545# => '0' & O"607",
    8#1546# => '1' & O"104",
    8#1547# => '0' & O"647",
    8#1550# => '1' & O"144",
    8#1551# => '0' & O"204",
    8#1552# => '1' & O"035",
    8#1553# => '0' & O"725",
    8#1554# => '0' & O"615",
    8#1555# => '1' & O"124",
    8#1556# => '0' & O"707",
    8#1557# => '1' & O"731",
    8#1560# => '0' & O"773",
    8#1561# => '1' & O"360",
    8#1562# => '0' & O"724",
    8#1563# => '0' & O"377",
    8#1564# => '0' & O"777",
    8#1565# => '0' & O"014",
    8#1566# => '1' & O"142",
    8#1567# => '1' & O"777",
    8#1570# => '0' & O"713",
    8#1571# => '1' & O"035",
    8#1572# => '0' & O"725",
    8#1573# => '1' & O"020",
    8#1574# => '0' & O"000",
    8#1575# => '0' & O"000",
    8#1576# => '1' & O"656",
    8#1577# => '1' & O"235",
    8#1600# => '0' & O"704",
    8#1601# => '1' & O"025",
    8#1602# => '1' & O"725",
    8#1603# => '1' & O"533",
    8#1604# => '0' & O"376",
    8#1605# => '1' & O"244",
    8#1606# => '1' & O"043",
    8#1607# => '1' & O"316",
    8#1610# => '0' & O"636",
    8#1611# => '1' & O"044",
    8#1612# => '1' & O"123",
    8#1613# => '0' & O"772",
    8#1614# => '1' & O"004",
    8#1615# => '0' & O"524",
    8#1616# => '1' & O"113",
    8#1617# => '0' & O"752",
    8#1620# => '1' & O"057",
    8#1621# => '0' & O"050",
    8#1622# => '0' & O"024",
    8#1623# => '1' & O"063",
    8#1624# => '0' & O"044",
    8#1625# => '0' & O"034",
    8#1626# => '1' & O"454",
    8#1627# => '1' & O"127",
    8#1630# => '1' & O"050",
    8#1631# => '1' & O"024",
    8#1632# => '1' & O"107",
    8#1633# => '0' & O"416",
    8#1634# => '0' & O"544",
    8#1635# => '1' & O"224",
    8#1636# => '0' & O"177",
    8#1637# => '1' & O"020",
    8#1640# => '0' & O"000",
    8#1641# => '0' & O"322",
    8#1642# => '0' & O"562",
    8#1643# => '0' & O"332",
    8#1644# => '1' & O"612",
    8#1645# => '1' & O"237",
    8#1646# => '0' & O"316",
    8#1647# => '0' & O"064",
    8#1650# => '0' & O"616",
    8#1651# => '1' & O"414",
    8#1652# => '0' & O"452",
    8#1653# => '0' & O"612",
    8#1654# => '0' & O"672",
    8#1655# => '1' & O"307",
    8#1656# => '0' & O"252",
    8#1657# => '0' & O"572",
    8#1660# => '1' & O"207",
    8#1661# => '1' & O"652",
    8#1662# => '0' & O"424",
    8#1663# => '0' & O"047",
    8#1664# => '1' & O"452",
    8#1665# => '0' & O"052",
    8#1666# => '1' & O"025",
    8#1667# => '1' & O"454",
    8#1670# => '1' & O"037",
    8#1671# => '0' & O"412",
    8#1672# => '1' & O"373",
    8#1673# => '0' & O"404",
    8#1674# => '1' & O"324",
    8#1675# => '0' & O"163",
    8#1676# => '1' & O"316",
    8#1677# => '1' & O"662",
    8#1700# => '1' & O"433",
    8#1701# => '1' & O"316",
    8#1702# => '0' & O"424",
    8#1703# => '1' & O"023",
    8#1704# => '1' & O"662",
    8#1705# => '0' & O"372",
    8#1706# => '0' & O"616",
    8#1707# => '0' & O"672",
    8#1710# => '1' & O"457",
    8#1711# => '0' & O"332",
    8#1712# => '0' & O"252",
    8#1713# => '1' & O"514",
    8#1714# => '0' & O"426",
    8#1715# => '0' & O"552",
    8#1716# => '1' & O"176",
    8#1717# => '1' & O"663",
    8#1720# => '1' & O"166",
    8#1721# => '1' & O"463",
    8#1722# => '0' & O"312",
    8#1723# => '1' & O"025",
    8#1724# => '1' & O"326",
    8#1725# => '0' & O"636",
    8#1726# => '1' & O"454",
    8#1727# => '1' & O"577",
    8#1730# => '0' & O"216",
    8#1731# => '0' & O"756",
    8#1732# => '0' & O"114",
    8#1733# => '0' & O"422",
    8#1734# => '0' & O"074",
    8#1735# => '0' & O"642",
    8#1736# => '1' & O"557",
    8#1737# => '1' & O"656",
    8#1740# => '0' & O"354",
    8#1741# => '1' & O"627",
    8#1742# => '0' & O"312",
    8#1743# => '0' & O"604",
    8#1744# => '1' & O"433",
    8#1745# => '0' & O"624",
    8#1746# => '1' & O"643",
    8#1747# => '0' & O"034",
    8#1750# => '1' & O"222",
    8#1751# => '1' & O"431",
    8#1752# => '0' & O"034",
    8#1753# => '0' & O"752",
    8#1754# => '0' & O"002",
    8#1755# => '1' & O"653",
    8#1756# => '1' & O"304",
    8#1757# => '1' & O"326",
    8#1760# => '1' & O"646",
    8#1761# => '0' & O"424",
    8#1762# => '1' & O"517",
    8#1763# => '1' & O"245",
    8#1764# => '1' & O"007",
    8#1765# => '1' & O"366",
    8#1766# => '0' & O"724",
    8#1767# => '1' & O"747",
    8#1770# => '0' & O"450",
    8#1771# => '0' & O"704",
    8#1772# => '0' & O"316",
    8#1773# => '0' & O"556",
    8#1774# => '0' & O"276",
    8#1775# => '0' & O"776",
    8#1776# => '1' & O"056",
    8#1777# => '0' & O"060",
    8#2000# => '0' & O"000",
    8#2001# => '1' & O"023",
    8#2002# => '0' & O"563",
    8#2003# => '1' & O"443",
    8#2004# => '0' & O"543",
    8#2005# => '1' & O"420",
    8#2006# => '0' & O"605",
    8#2007# => '0' & O"553",
    8#2010# => '1' & O"143",
    8#2011# => '0' & O"413",
    8#2012# => '1' & O"044",
    8#2013# => '0' & O"103",
    8#2014# => '0' & O"203",
    8#2015# => '0' & O"020",
    8#2016# => '0' & O"605",
    8#2017# => '1' & O"777",
    8#2020# => '0' & O"605",
    8#2021# => '0' & O"067",
    8#2022# => '1' & O"013",
    8#2023# => '1' & O"013",
    8#2024# => '1' & O"013",
    8#2025# => '1' & O"220",
    8#2026# => '0' & O"000",
    8#2027# => '0' & O"643",
    8#2030# => '1' & O"327",
    8#2031# => '0' & O"000",
    8#2032# => '1' & O"013",
    8#2033# => '1' & O"013",
    8#2034# => '1' & O"013",
    8#2035# => '0' & O"000",
    8#2036# => '0' & O"000",
    8#2037# => '0' & O"673",
    8#2040# => '0' & O"601",
    8#2041# => '1' & O"220",
    8#2042# => '1' & O"503",
    8#2043# => '0' & O"713",
    8#2044# => '0' & O"707",
    8#2045# => '0' & O"000",
    8#2046# => '0' & O"717",
    8#2047# => '0' & O"504",
    8#2050# => '0' & O"571",
    8#2051# => '0' & O"407",
    8#2052# => '0' & O"457",
    8#2053# => '0' & O"237",
    8#2054# => '1' & O"117",
    8#2055# => '1' & O"243",
    8#2056# => '0' & O"605",
    8#2057# => '0' & O"407",
    8#2060# => '0' & O"000",
    8#2061# => '0' & O"000",
    8#2062# => '1' & O"756",
    8#2063# => '1' & O"756",
    8#2064# => '0' & O"703",
    8#2065# => '1' & O"220",
    8#2066# => '0' & O"000",
    8#2067# => '0' & O"657",
    8#2070# => '0' & O"605",
    8#2071# => '1' & O"727",
    8#2072# => '1' & O"756",
    8#2073# => '0' & O"377",
    8#2074# => '0' & O"000",
    8#2075# => '0' & O"000",
    8#2076# => '1' & O"556",
    8#2077# => '0' & O"014",
    8#2100# => '0' & O"473",
    8#2101# => '0' & O"620",
    8#2102# => '0' & O"601",
    8#2103# => '1' & O"044",
    8#2104# => '1' & O"450",
    8#2105# => '0' & O"450",
    8#2106# => '0' & O"552",
    8#2107# => '0' & O"552",
    8#2110# => '1' & O"024",
    8#2111# => '1' & O"217",
    8#2112# => '1' & O"207",
    8#2113# => '0' & O"571",
    8#2114# => '0' & O"620",
    8#2115# => '0' & O"620",
    8#2116# => '0' & O"416",
    8#2117# => '0' & O"074",
    8#2120# => '1' & O"554",
    8#2121# => '0' & O"473",
    8#2122# => '0' & O"250",
    8#2123# => '1' & O"642",
    8#2124# => '0' & O"250",
    8#2125# => '0' & O"620",
    8#2126# => '0' & O"000",
    8#2127# => '0' & O"000",
    8#2130# => '0' & O"504",
    8#2131# => '0' & O"620",
    8#2132# => '1' & O"035",
    8#2133# => '0' & O"620",
    8#2134# => '1' & O"244",
    8#2135# => '0' & O"620",
    8#2136# => '0' & O"104",
    8#2137# => '0' & O"607",
    8#2140# => '0' & O"304",
    8#2141# => '1' & O"204",
    8#2142# => '1' & O"420",
    8#2143# => '1' & O"420",
    8#2144# => '1' & O"420",
    8#2145# => '1' & O"204",
    8#2146# => '0' & O"304",
    8#2147# => '0' & O"617",
    8#2150# => '0' & O"604",
    8#2151# => '0' & O"404",
    8#2152# => '0' & O"727",
    8#2153# => '0' & O"644",
    8#2154# => '0' & O"404",
    8#2155# => '0' & O"727",
    8#2156# => '0' & O"604",
    8#2157# => '0' & O"723",
    8#2160# => '1' & O"756",
    8#2161# => '1' & O"420",
    8#2162# => '1' & O"420",
    8#2163# => '0' & O"644",
    8#2164# => '0' & O"444",
    8#2165# => '0' & O"224",
    8#2166# => '0' & O"777",
    8#2167# => '1' & O"244",
    8#2170# => '0' & O"620",
    8#2171# => '1' & O"244",
    8#2172# => '1' & O"220",
    8#2173# => '0' & O"000",
    8#2174# => '1' & O"057",
    8#2175# => '0' & O"000",
    8#2176# => '0' & O"620",
    8#2177# => '0' & O"605",
    8#2200# => '0' & O"650",
    8#2201# => '0' & O"747",
    8#2202# => '1' & O"244",
    8#2203# => '1' & O"027",
    8#2204# => '1' & O"204",
    8#2205# => '1' & O"144",
    8#2206# => '0' & O"620",
    8#2207# => '0' & O"650",
    8#2210# => '0' & O"450",
    8#2211# => '1' & O"656",
    8#2212# => '0' & O"060",
    8#2213# => '1' & O"124",
    8#2214# => '1' & O"103",
    8#2215# => '0' & O"601",
    8#2216# => '1' & O"656",
    8#2217# => '0' & O"747",
    8#2220# => '0' & O"625",
    8#2221# => '1' & O"360",
    8#2222# => '1' & O"073",
    8#2223# => '0' & O"571",
    8#2224# => '0' & O"650",
    8#2225# => '0' & O"304",
    8#2226# => '1' & O"244",
    8#2227# => '0' & O"467",
    8#2230# => '0' & O"601",
    8#2231# => '1' & O"450",
    8#2232# => '0' & O"450",
    8#2233# => '1' & O"231",
    8#2234# => '0' & O"423",
    8#2235# => '0' & O"000",
    8#2236# => '0' & O"000",
    8#2237# => '1' & O"220",
    8#2240# => '0' & O"320",
    8#2241# => '0' & O"344",
    8#2242# => '1' & O"227",
    8#2243# => '0' & O"344",
    8#2244# => '0' & O"220",
    8#2245# => '0' & O"220",
    8#2246# => '0' & O"376",
    8#2247# => '0' & O"020",
    8#2250# => '0' & O"571",
    8#2251# => '0' & O"304",
    8#2252# => '0' & O"444",
    8#2253# => '0' & O"676",
    8#2254# => '1' & O"273",
    8#2255# => '0' & O"404",
    8#2256# => '1' & O"450",
    8#2257# => '1' & O"041",
    8#2260# => '1' & O"146",
    8#2261# => '0' & O"327",
    8#2262# => '0' & O"322",
    8#2263# => '0' & O"742",
    8#2264# => '0' & O"325",
    8#2265# => '0' & O"144",
    8#2266# => '1' & O"035",
    8#2267# => '0' & O"616",
    8#2270# => '1' & O"221",
    8#2271# => '1' & O"360",
    8#2272# => '1' & O"455",
    8#2273# => '0' & O"621",
    8#2274# => '1' & O"221",
    8#2275# => '1' & O"370",
    8#2276# => '1' & O"235",
    8#2277# => '1' & O"572",
    8#2300# => '1' & O"572",
    8#2301# => '1' & O"572",
    8#2302# => '1' & O"427",
    8#2303# => '0' & O"572",
    8#2304# => '1' & O"705",
    8#2305# => '0' & O"616",
    8#2306# => '0' & O"405",
    8#2307# => '1' & O"707",
    8#2310# => '0' & O"605",
    8#2311# => '0' & O"204",
    8#2312# => '0' & O"027",
    8#2313# => '0' & O"316",
    8#2314# => '1' & O"160",
    8#2315# => '0' & O"000",
    8#2316# => '1' & O"370",
    8#2317# => '0' & O"060",
    8#2320# => '1' & O"124",
    8#2321# => '1' & O"517",
    8#2322# => '1' & O"177",
    8#2323# => '0' & O"601",
    8#2324# => '0' & O"127",
    8#2325# => '0' & O"000",
    8#2326# => '0' & O"000",
    8#2327# => '0' & O"000",
    8#2330# => '0' & O"000",
    8#2331# => '0' & O"000",
    8#2332# => '0' & O"000",
    8#2333# => '0' & O"000",
    8#2334# => '0' & O"000",
    8#2335# => '0' & O"000",
    8#2336# => '0' & O"000",
    8#2337# => '0' & O"000",
    8#2340# => '0' & O"000",
    8#2341# => '0' & O"000",
    8#2342# => '0' & O"000",
    8#2343# => '0' & O"000",
    8#2344# => '0' & O"000",
    8#2345# => '0' & O"000",
    8#2346# => '0' & O"000",
    8#2347# => '0' & O"000",
    8#2350# => '0' & O"000",
    8#2351# => '0' & O"000",
    8#2352# => '0' & O"000",
    8#2353# => '0' & O"000",
    8#2354# => '0' & O"000",
    8#2355# => '0' & O"000",
    8#2356# => '0' & O"000",
    8#2357# => '0' & O"000",
    8#2360# => '0' & O"000",
    8#2361# => '0' & O"020",
    8#2362# => '0' & O"000",
    8#2363# => '0' & O"000",
    8#2364# => '0' & O"000",
    8#2365# => '1' & O"220",
    8#2366# => '0' & O"000",
    8#2367# => '0' & O"000",
    8#2370# => '0' & O"000",
    8#2371# => '0' & O"000",
    8#2372# => '0' & O"000",
    8#2373# => '0' & O"000",
    8#2374# => '0' & O"000",
    8#2375# => '0' & O"000",
    8#2376# => '0' & O"060",
    8#2377# => '1' & O"420",
    8#2400# => '1' & O"420",
    8#2401# => '0' & O"742",
    8#2402# => '0' & O"742",
    8#2403# => '0' & O"742",
    8#2404# => '0' & O"742",
    8#2405# => '0' & O"742",
    8#2406# => '0' & O"516",
    8#2407# => '1' & O"160",
    8#2410# => '0' & O"000",
    8#2411# => '1' & O"370",
    8#2412# => '0' & O"424",
    8#2413# => '1' & O"777",
    8#2414# => '1' & O"656",
    8#2415# => '1' & O"024",
    8#2416# => '1' & O"237",
    8#2417# => '1' & O"233",
    8#2420# => '0' & O"620",
    8#2421# => '0' & O"000",
    8#2422# => '0' & O"000",
    8#2423# => '0' & O"000",
    8#2424# => '0' & O"000",
    8#2425# => '1' & O"623",
    8#2426# => '0' & O"404",
    8#2427# => '1' & O"244",
    8#2430# => '1' & O"221",
    8#2431# => '0' & O"011",
    8#2432# => '1' & O"355",
    8#2433# => '0' & O"265",
    8#2434# => '0' & O"616",
    8#2435# => '0' & O"015",
    8#2436# => '0' & O"217",
    8#2437# => '0' & O"000",
    8#2440# => '0' & O"000",
    8#2441# => '0' & O"000",
    8#2442# => '0' & O"413",
    8#2443# => '1' & O"355",
    8#2444# => '0' & O"311",
    8#2445# => '0' & O"021",
    8#2446# => '1' & O"355",
    8#2447# => '0' & O"316",
    8#2450# => '0' & O"742",
    8#2451# => '0' & O"616",
    8#2452# => '0' & O"005",
    8#2453# => '1' & O"355",
    8#2454# => '0' & O"103",
    8#2455# => '0' & O"316",
    8#2456# => '1' & O"160",
    8#2457# => '0' & O"000",
    8#2460# => '1' & O"370",
    8#2461# => '0' & O"060",
    8#2462# => '1' & O"450",
    8#2463# => '0' & O"450",
    8#2464# => '0' & O"616",
    8#2465# => '0' & O"060",
    8#2466# => '1' & O"044",
    8#2467# => '1' & O"144",
    8#2470# => '1' & O"225",
    8#2471# => '0' & O"000",
    8#2472# => '0' & O"000",
    8#2473# => '0' & O"000",
    8#2474# => '0' & O"000",
    8#2475# => '0' & O"000",
    8#2476# => '0' & O"000",
    8#2477# => '0' & O"000",
    8#2500# => '0' & O"000",
    8#2501# => '0' & O"620",
    8#2502# => '1' & O"244",
    8#2503# => '0' & O"444",
    8#2504# => '0' & O"015",
    8#2505# => '0' & O"616",
    8#2506# => '1' & O"221",
    8#2507# => '0' & O"005",
    8#2510# => '0' & O"176",
    8#2511# => '0' & O"003",
    8#2512# => '1' & O"225",
    8#2513# => '0' & O"011",
    8#2514# => '1' & O"656",
    8#2515# => '1' & O"231",
    8#2516# => '0' & O"450",
    8#2517# => '0' & O"005",
    8#2520# => '1' & O"656",
    8#2521# => '0' & O"316",
    8#2522# => '0' & O"742",
    8#2523# => '1' & O"231",
    8#2524# => '0' & O"650",
    8#2525# => '1' & O"225",
    8#2526# => '0' & O"405",
    8#2527# => '0' & O"450",
    8#2530# => '0' & O"015",
    8#2531# => '0' & O"616",
    8#2532# => '0' & O"005",
    8#2533# => '1' & O"205",
    8#2534# => '0' & O"444",
    8#2535# => '0' & O"724",
    8#2536# => '0' & O"603",
    8#2537# => '0' & O"450",
    8#2540# => '0' & O"616",
    8#2541# => '0' & O"021",
    8#2542# => '0' & O"450",
    8#2543# => '0' & O"616",
    8#2544# => '0' & O"015",
    8#2545# => '0' & O"773",
    8#2546# => '0' & O"000",
    8#2547# => '0' & O"000",
    8#2550# => '0' & O"000",
    8#2551# => '0' & O"000",
    8#2552# => '0' & O"000",
    8#2553# => '0' & O"000",
    8#2554# => '0' & O"000",
    8#2555# => '0' & O"000",
    8#2556# => '0' & O"000",
    8#2557# => '0' & O"000",
    8#2560# => '0' & O"000",
    8#2561# => '0' & O"000",
    8#2562# => '0' & O"000",
    8#2563# => '0' & O"000",
    8#2564# => '0' & O"000",
    8#2565# => '1' & O"355",
    8#2566# => '1' & O"656",
    8#2567# => '0' & O"620",
    8#2570# => '0' & O"000",
    8#2571# => '0' & O"000",
    8#2572# => '0' & O"000",
    8#2573# => '1' & O"561",
    8#2574# => '1' & O"124",
    8#2575# => '0' & O"727",
    8#2576# => '0' & O"620",
    8#2577# => '0' & O"000",
    8#2600# => '0' & O"000",
    8#2601# => '0' & O"000",
    8#2602# => '0' & O"000",
    8#2603# => '0' & O"000",
    8#2604# => '0' & O"000",
    8#2605# => '0' & O"000",
    8#2606# => '0' & O"000",
    8#2607# => '0' & O"000",
    8#2610# => '0' & O"000",
    8#2611# => '0' & O"000",
    8#2612# => '0' & O"000",
    8#2613# => '0' & O"000",
    8#2614# => '0' & O"000",
    8#2615# => '0' & O"000",
    8#2616# => '0' & O"000",
    8#2617# => '0' & O"000",
    8#2620# => '0' & O"000",
    8#2621# => '0' & O"000",
    8#2622# => '0' & O"000",
    8#2623# => '0' & O"000",
    8#2624# => '0' & O"000",
    8#2625# => '0' & O"000",
    8#2626# => '0' & O"000",
    8#2627# => '0' & O"000",
    8#2630# => '0' & O"000",
    8#2631# => '0' & O"000",
    8#2632# => '0' & O"000",
    8#2633# => '0' & O"000",
    8#2634# => '0' & O"000",
    8#2635# => '0' & O"000",
    8#2636# => '0' & O"000",
    8#2637# => '0' & O"000",
    8#2640# => '0' & O"563",
    8#2641# => '0' & O"344",
    8#2642# => '1' & O"227",
    8#2643# => '0' & O"344",
    8#2644# => '0' & O"220",
    8#2645# => '0' & O"220",
    8#2646# => '0' & O"376",
    8#2647# => '0' & O"020",
    8#2650# => '0' & O"000",
    8#2651# => '0' & O"000",
    8#2652# => '0' & O"000",
    8#2653# => '0' & O"000",
    8#2654# => '0' & O"000",
    8#2655# => '0' & O"000",
    8#2656# => '0' & O"000",
    8#2657# => '0' & O"000",
    8#2660# => '0' & O"322",
    8#2661# => '0' & O"562",
    8#2662# => '0' & O"332",
    8#2663# => '0' & O"420",
    8#2664# => '1' & O"303",
    8#2665# => '0' & O"322",
    8#2666# => '0' & O"562",
    8#2667# => '0' & O"332",
    8#2670# => '1' & O"612",
    8#2671# => '1' & O"357",
    8#2672# => '0' & O"316",
    8#2673# => '0' & O"616",
    8#2674# => '1' & O"414",
    8#2675# => '0' & O"452",
    8#2676# => '0' & O"612",
    8#2677# => '0' & O"672",
    8#2700# => '1' & O"423",
    8#2701# => '0' & O"252",
    8#2702# => '0' & O"572",
    8#2703# => '1' & O"327",
    8#2704# => '1' & O"666",
    8#2705# => '1' & O"370",
    8#2706# => '1' & O"656",
    8#2707# => '1' & O"360",
    8#2710# => '0' & O"060",
    8#2711# => '0' & O"000",
    8#2712# => '0' & O"000",
    8#2713# => '0' & O"000",
    8#2714# => '0' & O"000",
    8#2715# => '0' & O"000",
    8#2716# => '0' & O"000",
    8#2717# => '0' & O"000",
    8#2720# => '0' & O"000",
    8#2721# => '0' & O"000",
    8#2722# => '0' & O"000",
    8#2723# => '0' & O"000",
    8#2724# => '0' & O"000",
    8#2725# => '0' & O"000",
    8#2726# => '0' & O"000",
    8#2727# => '0' & O"000",
    8#2730# => '0' & O"000",
    8#2731# => '0' & O"000",
    8#2732# => '0' & O"000",
    8#2733# => '0' & O"000",
    8#2734# => '0' & O"424",
    8#2735# => '1' & O"607",
    8#2736# => '0' & O"624",
    8#2737# => '1' & O"233",
    8#2740# => '1' & O"237",
    8#2741# => '0' & O"624",
    8#2742# => '1' & O"227",
    8#2743# => '1' & O"223",
    8#2744# => '0' & O"316",
    8#2745# => '0' & O"576",
    8#2746# => '0' & O"214",
    8#2747# => '0' & O"230",
    8#2750# => '0' & O"250",
    8#2751# => '0' & O"316",
    8#2752# => '1' & O"356",
    8#2753# => '1' & O"414",
    8#2754# => '0' & O"542",
    8#2755# => '1' & O"160",
    8#2756# => '1' & O"656",
    8#2757# => '0' & O"450",
    8#2760# => '1' & O"360",
    8#2761# => '1' & O"656",
    8#2762# => '0' & O"742",
    8#2763# => '0' & O"742",
    8#2764# => '1' & O"663",
    8#2765# => '0' & O"773",
    8#2766# => '0' & O"316",
    8#2767# => '0' & O"630",
    8#2770# => '1' & O"653",
    8#2771# => '0' & O"000",
    8#2772# => '0' & O"000",
    8#2773# => '0' & O"000",
    8#2774# => '0' & O"000",
    8#2775# => '0' & O"000",
    8#2776# => '0' & O"000",
    8#2777# => '0' & O"060",
    8#3000# => '1' & O"363",
    8#3001# => '0' & O"037",
    8#3002# => '0' & O"064",
    8#3003# => '0' & O"777",
    8#3004# => '0' & O"772",
    8#3005# => '0' & O"771",
    8#3006# => '1' & O"721",
    8#3007# => '0' & O"316",
    8#3010# => '0' & O"064",
    8#3011# => '0' & O"504",
    8#3012# => '0' & O"616",
    8#3013# => '1' & O"250",
    8#3014# => '1' & O"656",
    8#3015# => '0' & O"147",
    8#3016# => '1' & O"326",
    8#3017# => '1' & O"752",
    8#3020# => '0' & O"073",
    8#3021# => '1' & O"514",
    8#3022# => '1' & O"472",
    8#3023# => '0' & O"472",
    8#3024# => '0' & O"034",
    8#3025# => '0' & O"254",
    8#3026# => '0' & O"267",
    8#3027# => '1' & O"356",
    8#3030# => '1' & O"552",
    8#3031# => '0' & O"056",
    8#3032# => '1' & O"004",
    8#3033# => '0' & O"114",
    8#3034# => '0' & O"472",
    8#3035# => '0' & O"606",
    8#3036# => '0' & O"426",
    8#3037# => '1' & O"142",
    8#3040# => '0' & O"107",
    8#3041# => '1' & O"044",
    8#3042# => '1' & O"614",
    8#3043# => '0' & O"612",
    8#3044# => '0' & O"172",
    8#3045# => '0' & O"073",
    8#3046# => '0' & O"034",
    8#3047# => '0' & O"254",
    8#3050# => '0' & O"253",
    8#3051# => '0' & O"137",
    8#3052# => '1' & O"552",
    8#3053# => '0' & O"233",
    8#3054# => '0' & O"113",
    8#3055# => '1' & O"572",
    8#3056# => '0' & O"123",
    8#3057# => '0' & O"442",
    8#3060# => '0' & O"034",
    8#3061# => '1' & O"362",
    8#3062# => '0' & O"612",
    8#3063# => '1' & O"626",
    8#3064# => '0' & O"353",
    8#3065# => '1' & O"326",
    8#3066# => '1' & O"776",
    8#3067# => '1' & O"752",
    8#3070# => '1' & O"024",
    8#3071# => '0' & O"357",
    8#3072# => '0' & O"074",
    8#3073# => '1' & O"326",
    8#3074# => '0' & O"066",
    8#3075# => '1' & O"572",
    8#3076# => '1' & O"172",
    8#3077# => '0' & O"407",
    8#3100# => '0' & O"137",
    8#3101# => '1' & O"772",
    8#3102# => '1' & O"456",
    8#3103# => '1' & O"742",
    8#3104# => '1' & O"742",
    8#3105# => '0' & O"426",
    8#3106# => '1' & O"572",
    8#3107# => '0' & O"427",
    8#3110# => '1' & O"362",
    8#3111# => '1' & O"562",
    8#3112# => '1' & O"326",
    8#3113# => '1' & O"456",
    8#3114# => '1' & O"024",
    8#3115# => '0' & O"527",
    8#3116# => '1' & O"652",
    8#3117# => '0' & O"052",
    8#3120# => '0' & O"672",
    8#3121# => '0' & O"523",
    8#3122# => '0' & O"252",
    8#3123# => '0' & O"572",
    8#3124# => '1' & O"652",
    8#3125# => '0' & O"524",
    8#3126# => '1' & O"773",
    8#3127# => '1' & O"003",
    8#3130# => '0' & O"000",
    8#3131# => '0' & O"000",
    8#3132# => '0' & O"000",
    8#3133# => '0' & O"000",
    8#3134# => '0' & O"000",
    8#3135# => '0' & O"000",
    8#3136# => '0' & O"000",
    8#3137# => '0' & O"000",
    8#3140# => '0' & O"000",
    8#3141# => '0' & O"000",
    8#3142# => '0' & O"000",
    8#3143# => '1' & O"323",
    8#3144# => '1' & O"223",
    8#3145# => '0' & O"616",
    8#3146# => '0' & O"316",
    8#3147# => '0' & O"542",
    8#3150# => '1' & O"160",
    8#3151# => '1' & O"656",
    8#3152# => '0' & O"616",
    8#3153# => '1' & O"757",
    8#3154# => '0' & O"000",
    8#3155# => '0' & O"000",
    8#3156# => '0' & O"000",
    8#3157# => '0' & O"000",
    8#3160# => '0' & O"000",
    8#3161# => '0' & O"000",
    8#3162# => '1' & O"007",
    8#3163# => '0' & O"731",
    8#3164# => '0' & O"064",
    8#3165# => '0' & O"220",
    8#3166# => '0' & O"724",
    8#3167# => '0' & O"747",
    8#3170# => '0' & O"450",
    8#3171# => '0' & O"316",
    8#3172# => '0' & O"060",
    8#3173# => '0' & O"000",
    8#3174# => '1' & O"244",
    8#3175# => '0' & O"621",
    8#3176# => '0' & O"620",
    8#3177# => '0' & O"145",
    8#3200# => '0' & O"620",
    8#3201# => '0' & O"416",
    8#3202# => '0' & O"416",
    8#3203# => '0' & O"731",
    8#3204# => '1' & O"572",
    8#3205# => '1' & O"037",
    8#3206# => '0' & O"763",
    8#3207# => '1' & O"572",
    8#3210# => '1' & O"067",
    8#3211# => '0' & O"230",
    8#3212# => '0' & O"530",
    8#3213# => '0' & O"430",
    8#3214# => '0' & O"773",
    8#3215# => '1' & O"572",
    8#3216# => '1' & O"147",
    8#3217# => '0' & O"430",
    8#3220# => '0' & O"530",
    8#3221# => '0' & O"330",
    8#3222# => '0' & O"530",
    8#3223# => '1' & O"130",
    8#3224# => '0' & O"230",
    8#3225# => '0' & O"330",
    8#3226# => '0' & O"730",
    8#3227# => '0' & O"552",
    8#3230# => '0' & O"771",
    8#3231# => '0' & O"330",
    8#3232# => '0' & O"730",
    8#3233# => '1' & O"030",
    8#3234# => '0' & O"530",
    8#3235# => '0' & O"430",
    8#3236# => '0' & O"130",
    8#3237# => '0' & O"130",
    8#3240# => '0' & O"730",
    8#3241# => '1' & O"030",
    8#3242# => '0' & O"430",
    8#3243# => '0' & O"773",
    8#3244# => '0' & O"014",
    8#3245# => '0' & O"416",
    8#3246# => '0' & O"074",
    8#3247# => '1' & O"454",
    8#3250# => '1' & O"227",
    8#3251# => '1' & O"376",
    8#3252# => '1' & O"656",
    8#3253# => '1' & O"160",
    8#3254# => '0' & O"244",
    8#3255# => '1' & O"370",
    8#3256# => '1' & O"656",
    8#3257# => '1' & O"344",
    8#3260# => '0' & O"056",
    8#3261# => '0' & O"124",
    8#3262# => '1' & O"757",
    8#3263# => '0' & O"627",
    8#3264# => '0' & O"456",
    8#3265# => '1' & O"656",
    8#3266# => '0' & O"316",
    8#3267# => '1' & O"160",
    8#3270# => '0' & O"216",
    8#3271# => '1' & O"656",
    8#3272# => '1' & O"360",
    8#3273# => '0' & O"623",
    8#3274# => '0' & O"176",
    8#3275# => '0' & O"037",
    8#3276# => '0' & O"172",
    8#3277# => '0' & O"037",
    8#3300# => '0' & O"152",
    8#3301# => '1' & O"423",
    8#3302# => '0' & O"034",
    8#3303# => '1' & O"457",
    8#3304# => '0' & O"034",
    8#3305# => '0' & O"354",
    8#3306# => '1' & O"443",
    8#3307# => '0' & O"023",
    8#3310# => '0' & O"552",
    8#3311# => '1' & O"401",
    8#3312# => '0' & O"420",
    8#3313# => '0' & O"162",
    8#3314# => '0' & O"037",
    8#3315# => '1' & O"652",
    8#3316# => '1' & O"314",
    8#3317# => '0' & O"652",
    8#3320# => '1' & O"527",
    8#3321# => '0' & O"552",
    8#3322# => '0' & O"152",
    8#3323# => '0' & O"023",
    8#3324# => '0' & O"416",
    8#3325# => '1' & O"656",
    8#3326# => '1' & O"356",
    8#3327# => '1' & O"742",
    8#3330# => '0' & O"256",
    8#3331# => '1' & O"453",
    8#3332# => '1' & O"656",
    8#3333# => '1' & O"116",
    8#3334# => '0' & O"776",
    8#3335# => '1' & O"414",
    8#3336# => '0' & O"466",
    8#3337# => '1' & O"716",
    8#3340# => '1' & O"577",
    8#3341# => '1' & O"516",
    8#3342# => '0' & O"416",
    8#3343# => '1' & O"716",
    8#3344# => '1' & O"617",
    8#3345# => '1' & O"776",
    8#3346# => '1' & O"456",
    8#3347# => '1' & O"731",
    8#3350# => '1' & O"314",
    8#3351# => '1' & O"731",
    8#3352# => '0' & O"216",
    8#3353# => '0' & O"062",
    8#3354# => '1' & O"216",
    8#3355# => '1' & O"456",
    8#3356# => '1' & O"626",
    8#3357# => '1' & O"567",
    8#3360# => '1' & O"656",
    8#3361# => '1' & O"052",
    8#3362# => '0' & O"752",
    8#3363# => '1' & O"451",
    8#3364# => '1' & O"044",
    8#3365# => '0' & O"420",
    8#3366# => '0' & O"002",
    8#3367# => '1' & O"753",
    8#3370# => '1' & O"222",
    8#3371# => '1' & O"752",
    8#3372# => '0' & O"060",
    8#3373# => '1' & O"224",
    8#3374# => '1' & O"773",
    8#3375# => '1' & O"020",
    8#3376# => '0' & O"620",
    8#3377# => '0' & O"000",
    8#3400# => '0' & O"027",
    8#3401# => '1' & O"213",
    8#3402# => '0' & O"027",
    8#3403# => '0' & O"027",
    8#3404# => '0' & O"027",
    8#3405# => '0' & O"067",
    8#3406# => '0' & O"027",
    8#3407# => '0' & O"107",
    8#3410# => '0' & O"027",
    8#3411# => '1' & O"237",
    8#3412# => '0' & O"027",
    8#3413# => '0' & O"027",
    8#3414# => '0' & O"027",
    8#3415# => '1' & O"223",
    8#3416# => '0' & O"027",
    8#3417# => '1' & O"130",
    8#3420# => '1' & O"117",
    8#3421# => '1' & O"227",
    8#3422# => '0' & O"303",
    8#3423# => '0' & O"177",
    8#3424# => '0' & O"430",
    8#3425# => '0' & O"767",
    8#3426# => '0' & O"027",
    8#3427# => '1' & O"030",
    8#3430# => '1' & O"117",
    8#3431# => '1' & O"243",
    8#3432# => '0' & O"753",
    8#3433# => '0' & O"763",
    8#3434# => '0' & O"130",
    8#3435# => '0' & O"767",
    8#3436# => '0' & O"027",
    8#3437# => '0' & O"530",
    8#3440# => '1' & O"117",
    8#3441# => '0' & O"237",
    8#3442# => '1' & O"103",
    8#3443# => '1' & O"507",
    8#3444# => '0' & O"030",
    8#3445# => '0' & O"767",
    8#3446# => '0' & O"027",
    8#3447# => '0' & O"047",
    8#3450# => '0' & O"027",
    8#3451# => '0' & O"267",
    8#3452# => '0' & O"027",
    8#3453# => '0' & O"027",
    8#3454# => '0' & O"027",
    8#3455# => '0' & O"277",
    8#3456# => '0' & O"027",
    8#3457# => '0' & O"337",
    8#3460# => '0' & O"630",
    8#3461# => '1' & O"117",
    8#3462# => '0' & O"077",
    8#3463# => '0' & O"137",
    8#3464# => '0' & O"730",
    8#3465# => '0' & O"767",
    8#3466# => '0' & O"027",
    8#3467# => '1' & O"767",
    8#3470# => '1' & O"356",
    8#3471# => '0' & O"065",
    8#3472# => '0' & O"723",
    8#3473# => '1' & O"073",
    8#3474# => '0' & O"713",
    8#3475# => '0' & O"620",
    8#3476# => '1' & O"124",
    8#3477# => '0' & O"367",
    8#3500# => '0' & O"064",
    8#3501# => '0' & O"176",
    8#3502# => '1' & O"773",
    8#3503# => '0' & O"552",
    8#3504# => '0' & O"552",
    8#3505# => '0' & O"672",
    8#3506# => '1' & O"773",
    8#3507# => '0' & O"447",
    8#3510# => '1' & O"106",
    8#3511# => '0' & O"752",
    8#3512# => '0' & O"443",
    8#3513# => '1' & O"656",
    8#3514# => '1' & O"250",
    8#3515# => '0' & O"130",
    8#3516# => '0' & O"330",
    8#3517# => '0' & O"106",
    8#3520# => '1' & O"773",
    8#3521# => '0' & O"630",
    8#3522# => '1' & O"214",
    8#3523# => '0' & O"102",
    8#3524# => '1' & O"773",
    8#3525# => '1' & O"014",
    8#3526# => '1' & O"322",
    8#3527# => '0' & O"714",
    8#3530# => '0' & O"630",
    8#3531# => '0' & O"714",
    8#3532# => '0' & O"102",
    8#3533# => '1' & O"773",
    8#3534# => '0' & O"250",
    8#3535# => '0' & O"514",
    8#3536# => '1' & O"322",
    8#3537# => '1' & O"322",
    8#3540# => '1' & O"322",
    8#3541# => '1' & O"322",
    8#3542# => '1' & O"456",
    8#3543# => '1' & O"562",
    8#3544# => '1' & O"352",
    8#3545# => '1' & O"014",
    8#3546# => '1' & O"542",
    8#3547# => '1' & O"314",
    8#3550# => '1' & O"742",
    8#3551# => '1' & O"742",
    8#3552# => '1' & O"576",
    8#3553# => '1' & O"456",
    8#3554# => '0' & O"044",
    8#3555# => '0' & O"245",
    8#3556# => '0' & O"245",
    8#3557# => '0' & O"024",
    8#3560# => '1' & O"063",
    8#3561# => '1' & O"233",
    8#3562# => '1' & O"204",
    8#3563# => '1' & O"223",
    8#3564# => '0' & O"012",
    8#3565# => '1' & O"043",
    8#3566# => '0' & O"052",
    8#3567# => '0' & O"037",
    8#3570# => '0' & O"000",
    8#3571# => '0' & O"000",
    8#3572# => '0' & O"330",
    8#3573# => '1' & O"117",
    8#3574# => '0' & O"230",
    8#3575# => '1' & O"117",
    8#3576# => '0' & O"620",
    8#3577# => '0' & O"024",
    8#3600# => '0' & O"007",
    8#3601# => '1' & O"024",
    8#3602# => '0' & O"663",
    8#3603# => '1' & O"050",
    8#3604# => '1' & O"044",
    8#3605# => '1' & O"414",
    8#3606# => '0' & O"316",
    8#3607# => '0' & O"320",
    8#3610# => '1' & O"452",
    8#3611# => '1' & O"552",
    8#3612# => '1' & O"452",
    8#3613# => '1' & O"227",
    8#3614# => '1' & O"004",
    8#3615# => '0' & O"207",
    8#3616# => '1' & O"224",
    8#3617# => '0' & O"713",
    8#3620# => '1' & O"244",
    8#3621# => '1' & O"160",
    8#3622# => '1' & O"133",
    8#3623# => '1' & O"160",
    8#3624# => '1' & O"224",
    8#3625# => '1' & O"157",
    8#3626# => '1' & O"656",
    8#3627# => '0' & O"616",
    8#3630# => '1' & O"106",
    8#3631# => '1' & O"360",
    8#3632# => '1' & O"233",
    8#3633# => '1' & O"370",
    8#3634# => '1' & O"414",
    8#3635# => '0' & O"642",
    8#3636# => '1' & O"203",
    8#3637# => '0' & O"316",
    8#3640# => '1' & O"656",
    8#3641# => '0' & O"426",
    8#3642# => '0' & O"265",
    8#3643# => '0' & O"275",
    8#3644# => '0' & O"275",
    8#3645# => '0' & O"275",
    8#3646# => '0' & O"275",
    8#3647# => '0' & O"335",
    8#3650# => '1' & O"250",
    8#3651# => '1' & O"050",
    8#3652# => '0' & O"050",
    8#3653# => '1' & O"224",
    8#3654# => '0' & O"777",
    8#3655# => '0' & O"114",
    8#3656# => '1' & O"762",
    8#3657# => '0' & O"777",
    8#3660# => '0' & O"614",
    8#3661# => '1' & O"742",
    8#3662# => '1' & O"213",
    8#3663# => '0' & O"714",
    8#3664# => '1' & O"742",
    8#3665# => '0' & O"102",
    8#3666# => '1' & O"343",
    8#3667# => '1' & O"217",
    8#3670# => '1' & O"362",
    8#3671# => '1' & O"114",
    8#3672# => '1' & O"742",
    8#3673# => '0' & O"067",
    8#3674# => '1' & O"214",
    8#3675# => '1' & O"742",
    8#3676# => '0' & O"102",
    8#3677# => '1' & O"407",
    8#3700# => '1' & O"227",
    8#3701# => '0' & O"322",
    8#3702# => '1' & O"362",
    8#3703# => '1' & O"314",
    8#3704# => '1' & O"742",
    8#3705# => '1' & O"453",
    8#3706# => '1' & O"356",
    8#3707# => '1' & O"414",
    8#3710# => '1' & O"742",
    8#3711# => '1' & O"237",
    8#3712# => '0' & O"106",
    8#3713# => '1' & O"467",
    8#3714# => '0' & O"047",
    8#3715# => '1' & O"356",
    8#3716# => '1' & O"314",
    8#3717# => '1' & O"742",
    8#3720# => '0' & O"147",
    8#3721# => '1' & O"250",
    8#3722# => '0' & O"322",
    8#3723# => '0' & O"214",
    8#3724# => '0' & O"012",
    8#3725# => '1' & O"543",
    8#3726# => '0' & O"430",
    8#3727# => '1' & O"547",
    8#3730# => '0' & O"630",
    8#3731# => '0' & O"250",
    8#3732# => '0' & O"316",
    8#3733# => '1' & O"414",
    8#3734# => '0' & O"056",
    8#3735# => '1' & O"160",
    8#3736# => '1' & O"056",
    8#3737# => '1' & O"370",
    8#3740# => '0' & O"142",
    8#3741# => '1' & O"623",
    8#3742# => '1' & O"655",
    8#3743# => '1' & O"360",
    8#3744# => '1' & O"056",
    8#3745# => '0' & O"742",
    8#3746# => '1' & O"567",
    8#3747# => '1' & O"306",
    8#3750# => '1' & O"656",
    8#3751# => '1' & O"655",
    8#3752# => '0' & O"773",
    8#3753# => '0' & O"662",
    8#3754# => '1' & O"767",
    8#3755# => '1' & O"656",
    8#3756# => '0' & O"416",
    8#3757# => '1' & O"014",
    8#3760# => '0' & O"422",
    8#3761# => '0' & O"614",
    8#3762# => '0' & O"422",
    8#3763# => '0' & O"422",
    8#3764# => '0' & O"422",
    8#3765# => '1' & O"414",
    8#3766# => '1' & O"752",
    8#3767# => '1' & O"142",
    8#3770# => '1' & O"763",
    8#3771# => '1' & O"552",
    8#3772# => '0' & O"406",
    8#3773# => '1' & O"737",
    8#3774# => '1' & O"656",
    8#3775# => '0' & O"060",
    8#3776# => '0' & O"316",
    8#3777# => '0' & O"455"
  );  -- End 45 ROM

  constant ROM_55 : RomType := (
    8#0000# => '0' & O"575",
    8#0001# => '1' & O"364",
    8#0002# => '0' & O"477",
    8#0003# => '0' & O"564",
    8#0004# => '0' & O"757",
    8#0005# => '0' & O"504",
    8#0006# => '1' & O"414",
    8#0007# => '0' & O"420",
    8#0010# => '0' & O"742",
    8#0011# => '1' & O"145",
    8#0012# => '1' & O"414",
    8#0013# => '0' & O"530",
    8#0014# => '0' & O"030",
    8#0015# => '1' & O"654",
    8#0016# => '0' & O"057",
    8#0017# => '1' & O"656",
    8#0020# => '0' & O"416",
    8#0021# => '1' & O"414",
    8#0022# => '0' & O"230",
    8#0023# => '0' & O"330",
    8#0024# => '1' & O"314",
    8#0025# => '0' & O"217",
    8#0026# => '0' & O"561",
    8#0027# => '0' & O"624",
    8#0030# => '0' & O"027",
    8#0031# => '0' & O"504",
    8#0032# => '1' & O"204",
    8#0033# => '1' & O"104",
    8#0034# => '1' & O"414",
    8#0035# => '0' & O"564",
    8#0036# => '0' & O"013",
    8#0037# => '0' & O"561",
    8#0040# => '0' & O"624",
    8#0041# => '0' & O"033",
    8#0042# => '0' & O"153",
    8#0043# => '0' & O"752",
    8#0044# => '1' & O"160",
    8#0045# => '1' & O"656",
    8#0046# => '1' & O"563",
    8#0047# => '0' & O"450",
    8#0050# => '0' & O"504",
    8#0051# => '1' & O"541",
    8#0052# => '0' & O"773",
    8#0053# => '0' & O"144",
    8#0054# => '0' & O"244",
    8#0055# => '1' & O"414",
    8#0056# => '0' & O"056",
    8#0057# => '1' & O"420",
    8#0060# => '0' & O"456",
    8#0061# => '1' & O"343",
    8#0062# => '1' & O"364",
    8#0063# => '0' & O"107",
    8#0064# => '0' & O"621",
    8#0065# => '0' & O"561",
    8#0066# => '0' & O"424",
    8#0067# => '1' & O"023",
    8#0070# => '0' & O"616",
    8#0071# => '0' & O"005",
    8#0072# => '1' & O"037",
    8#0073# => '0' & O"614",
    8#0074# => '0' & O"250",
    8#0075# => '0' & O"060",
    8#0076# => '0' & O"564",
    8#0077# => '0' & O"603",
    8#0100# => '0' & O"355",
    8#0101# => '1' & O"130",
    8#0102# => '1' & O"363",
    8#0103# => '0' & O"564",
    8#0104# => '0' & O"643",
    8#0105# => '0' & O"000",
    8#0106# => '0' & O"621",
    8#0107# => '0' & O"724",
    8#0110# => '0' & O"453",
    8#0111# => '0' & O"450",
    8#0112# => '1' & O"121",
    8#0113# => '1' & O"037",
    8#0114# => '0' & O"616",
    8#0115# => '0' & O"316",
    8#0116# => '1' & O"414",
    8#0117# => '0' & O"542",
    8#0120# => '0' & O"752",
    8#0121# => '1' & O"443",
    8#0122# => '0' & O"000",
    8#0123# => '0' & O"323",
    8#0124# => '1' & O"141",
    8#0125# => '1' & O"037",
    8#0126# => '0' & O"000",
    8#0127# => '0' & O"242",
    8#0130# => '0' & O"242",
    8#0131# => '1' & O"243",
    8#0132# => '0' & O"250",
    8#0133# => '1' & O"007",
    8#0134# => '0' & O"420",
    8#0135# => '1' & O"364",
    8#0136# => '0' & O"167",
    8#0137# => '1' & O"131",
    8#0140# => '0' & O"604",
    8#0141# => '1' & O"141",
    8#0142# => '1' & O"414",
    8#0143# => '0' & O"043",
    8#0144# => '1' & O"220",
    8#0145# => '0' & O"544",
    8#0146# => '0' & O"404",
    8#0147# => '0' & O"650",
    8#0150# => '1' & O"431",
    8#0151# => '0' & O"311",
    8#0152# => '0' & O"303",
    8#0153# => '0' & O"250",
    8#0154# => '0' & O"614",
    8#0155# => '0' & O"742",
    8#0156# => '0' & O"542",
    8#0157# => '0' & O"537",
    8#0160# => '0' & O"250",
    8#0161# => '1' & O"552",
    8#0162# => '1' & O"552",
    8#0163# => '1' & O"255",
    8#0164# => '1' & O"121",
    8#0165# => '0' & O"005",
    8#0166# => '0' & O"311",
    8#0167# => '0' & O"450",
    8#0170# => '0' & O"415",
    8#0171# => '0' & O"650",
    8#0172# => '0' & O"450",
    8#0173# => '1' & O"656",
    8#0174# => '1' & O"104",
    8#0175# => '0' & O"243",
    8#0176# => '0' & O"616",
    8#0177# => '0' & O"424",
    8#0200# => '0' & O"657",
    8#0201# => '1' & O"541",
    8#0202# => '0' & O"015",
    8#0203# => '1' & O"613",
    8#0204# => '0' & O"176",
    8#0205# => '1' & O"773",
    8#0206# => '0' & O"255",
    8#0207# => '0' & O"220",
    8#0210# => '0' & O"524",
    8#0211# => '1' & O"037",
    8#0212# => '1' & O"224",
    8#0213# => '0' & O"627",
    8#0214# => '1' & O"244",
    8#0215# => '0' & O"650",
    8#0216# => '0' & O"450",
    8#0217# => '0' & O"456",
    8#0220# => '1' & O"343",
    8#0221# => '0' & O"355",
    8#0222# => '0' & O"030",
    8#0223# => '1' & O"363",
    8#0224# => '0' & O"564",
    8#0225# => '1' & O"073",
    8#0226# => '0' & O"064",
    8#0227# => '1' & O"650",
    8#0230# => '0' & O"316",
    8#0231# => '0' & O"752",
    8#0232# => '1' & O"414",
    8#0233# => '0' & O"624",
    8#0234# => '1' & O"173",
    8#0235# => '0' & O"742",
    8#0236# => '1' & O"314",
    8#0237# => '1' & O"160",
    8#0240# => '1' & O"056",
    8#0241# => '1' & O"360",
    8#0242# => '0' & O"450",
    8#0243# => '1' & O"056",
    8#0244# => '0' & O"742",
    8#0245# => '1' & O"177",
    8#0246# => '0' & O"216",
    8#0247# => '0' & O"060",
    8#0250# => '0' & O"250",
    8#0251# => '0' & O"461",
    8#0252# => '0' & O"565",
    8#0253# => '1' & O"451",
    8#0254# => '0' & O"005",
    8#0255# => '0' & O"311",
    8#0256# => '1' & O"007",
    8#0257# => '0' & O"561",
    8#0260# => '0' & O"424",
    8#0261# => '1' & O"317",
    8#0262# => '0' & O"376",
    8#0263# => '0' & O"444",
    8#0264# => '0' & O"504",
    8#0265# => '1' & O"204",
    8#0266# => '0' & O"000",
    8#0267# => '1' & O"056",
    8#0270# => '1' & O"264",
    8#0271# => '0' & O"420",
    8#0272# => '0' & O"355",
    8#0273# => '0' & O"130",
    8#0274# => '0' & O"250",
    8#0275# => '0' & O"564",
    8#0276# => '0' & O"117",
    8#0277# => '0' & O"621",
    8#0300# => '0' & O"724",
    8#0301# => '1' & O"417",
    8#0302# => '0' & O"450",
    8#0303# => '1' & O"451",
    8#0304# => '1' & O"256",
    8#0305# => '1' & O"037",
    8#0306# => '1' & O"364",
    8#0307# => '1' & O"143",
    8#0310# => '0' & O"220",
    8#0311# => '0' & O"000",
    8#0312# => '0' & O"144",
    8#0313# => '1' & O"420",
    8#0314# => '1' & O"541",
    8#0315# => '1' & O"224",
    8#0316# => '1' & O"523",
    8#0317# => '1' & O"124",
    8#0320# => '0' & O"723",
    8#0321# => '1' & O"121",
    8#0322# => '0' & O"005",
    8#0323# => '0' & O"000",
    8#0324# => '0' & O"450",
    8#0325# => '1' & O"144",
    8#0326# => '0' & O"415",
    8#0327# => '1' & O"037",
    8#0330# => '0' & O"304",
    8#0331# => '1' & O"344",
    8#0332# => '1' & O"004",
    8#0333# => '0' & O"060",
    8#0334# => '1' & O"360",
    8#0335# => '1' & O"656",
    8#0336# => '0' & O"742",
    8#0337# => '0' & O"223",
    8#0340# => '1' & O"650",
    8#0341# => '1' & O"743",
    8#0342# => '0' & O"650",
    8#0343# => '0' & O"104",
    8#0344# => '1' & O"124",
    8#0345# => '1' & O"643",
    8#0346# => '0' & O"263",
    8#0347# => '1' & O"020",
    8#0350# => '1' & O"656",
    8#0351# => '0' & O"312",
    8#0352# => '0' & O"014",
    8#0353# => '0' & O"530",
    8#0354# => '0' & O"252",
    8#0355# => '1' & O"656",
    8#0356# => '0' & O"672",
    8#0357# => '0' & O"263",
    8#0360# => '0' & O"112",
    8#0361# => '1' & O"717",
    8#0362# => '0' & O"263",
    8#0363# => '0' & O"616",
    8#0364# => '0' & O"424",
    8#0365# => '1' & O"463",
    8#0366# => '0' & O"764",
    8#0367# => '1' & O"067",
    8#0370# => '1' & O"214",
    8#0371# => '0' & O"130",
    8#0372# => '0' & O"714",
    8#0373# => '0' & O"230",
    8#0374# => '0' & O"564",
    8#0375# => '0' & O"333",
    8#0376# => '0' & O"764",
    8#0377# => '1' & O"413",
    8#0400# => '0' & O"104",
    8#0401# => '0' & O"347",
    8#0402# => '0' & O"332",
    8#0403# => '1' & O"771",
    8#0404# => '0' & O"000",
    8#0405# => '0' & O"542",
    8#0406# => '1' & O"363",
    8#0407# => '0' & O"601",
    8#0410# => '1' & O"024",
    8#0411# => '1' & O"337",
    8#0412# => '0' & O"216",
    8#0413# => '1' & O"347",
    8#0414# => '0' & O"564",
    8#0415# => '1' & O"017",
    8#0416# => '1' & O"364",
    8#0417# => '0' & O"567",
    8#0420# => '0' & O"542",
    8#0421# => '0' & O"167",
    8#0422# => '0' & O"250",
    8#0423# => '0' & O"176",
    8#0424# => '0' & O"627",
    8#0425# => '0' & O"250",
    8#0426# => '0' & O"367",
    8#0427# => '0' & O"324",
    8#0430# => '0' & O"577",
    8#0431# => '1' & O"324",
    8#0432# => '1' & O"257",
    8#0433# => '1' & O"364",
    8#0434# => '1' & O"473",
    8#0435# => '0' & O"250",
    8#0436# => '0' & O"676",
    8#0437# => '0' & O"207",
    8#0440# => '1' & O"675",
    8#0441# => '0' & O"250",
    8#0442# => '0' & O"542",
    8#0443# => '0' & O"303",
    8#0444# => '1' & O"221",
    8#0445# => '0' & O"757",
    8#0446# => '0' & O"124",
    8#0447# => '0' & O"073",
    8#0450# => '1' & O"656",
    8#0451# => '0' & O"250",
    8#0452# => '1' & O"014",
    8#0453# => '0' & O"272",
    8#0454# => '1' & O"473",
    8#0455# => '0' & O"130",
    8#0456# => '1' & O"477",
    8#0457# => '0' & O"000",
    8#0460# => '0' & O"542",
    8#0461# => '0' & O"413",
    8#0462# => '1' & O"221",
    8#0463# => '1' & O"747",
    8#0464# => '0' & O"216",
    8#0465# => '1' & O"057",
    8#0466# => '1' & O"364",
    8#0467# => '0' & O"107",
    8#0470# => '0' & O"250",
    8#0471# => '0' & O"575",
    8#0472# => '1' & O"124",
    8#0473# => '0' & O"323",
    8#0474# => '1' & O"057",
    8#0475# => '1' & O"515",
    8#0476# => '0' & O"224",
    8#0477# => '0' & O"233",
    8#0500# => '0' & O"764",
    8#0501# => '1' & O"733",
    8#0502# => '0' & O"542",
    8#0503# => '0' & O"477",
    8#0504# => '1' & O"221",
    8#0505# => '1' & O"661",
    8#0506# => '1' & O"701",
    8#0507# => '0' & O"250",
    8#0510# => '0' & O"332",
    8#0511# => '0' & O"772",
    8#0512# => '0' & O"204",
    8#0513# => '0' & O"343",
    8#0514# => '0' & O"564",
    8#0515# => '0' & O"757",
    8#0516# => '1' & O"220",
    8#0517# => '0' & O"542",
    8#0520# => '1' & O"277",
    8#0521# => '1' & O"221",
    8#0522# => '0' & O"056",
    8#0523# => '1' & O"515",
    8#0524# => '0' & O"064",
    8#0525# => '0' & O"347",
    8#0526# => '0' & O"724",
    8#0527# => '0' & O"553",
    8#0530# => '1' & O"056",
    8#0531# => '0' & O"450",
    8#0532# => '1' & O"104",
    8#0533# => '0' & O"717",
    8#0534# => '0' & O"420",
    8#0535# => '0' & O"542",
    8#0536# => '0' & O"027",
    8#0537# => '1' & O"044",
    8#0540# => '0' & O"344",
    8#0541# => '1' & O"344",
    8#0542# => '0' & O"060",
    8#0543# => '0' & O"000",
    8#0544# => '1' & O"220",
    8#0545# => '0' & O"576",
    8#0546# => '0' & O"676",
    8#0547# => '1' & O"527",
    8#0550# => '1' & O"656",
    8#0551# => '0' & O"250",
    8#0552# => '0' & O"014",
    8#0553# => '0' & O"602",
    8#0554# => '1' & O"242",
    8#0555# => '1' & O"437",
    8#0556# => '1' & O"642",
    8#0557# => '0' & O"250",
    8#0560# => '1' & O"656",
    8#0561# => '1' & O"675",
    8#0562# => '0' & O"117",
    8#0563# => '0' & O"316",
    8#0564# => '1' & O"356",
    8#0565# => '1' & O"414",
    8#0566# => '0' & O"562",
    8#0567# => '0' & O"776",
    8#0570# => '0' & O"776",
    8#0571# => '1' & O"056",
    8#0572# => '1' & O"727",
    8#0573# => '0' & O"621",
    8#0574# => '0' & O"561",
    8#0575# => '1' & O"515",
    8#0576# => '0' & O"650",
    8#0577# => '1' & O"656",
    8#0600# => '0' & O"450",
    8#0601# => '0' & O"552",
    8#0602# => '0' & O"552",
    8#0603# => '0' & O"471",
    8#0604# => '1' & O"043",
    8#0605# => '0' & O"650",
    8#0606# => '0' & O"450",
    8#0607# => '0' & O"060",
    8#0610# => '0' & O"064",
    8#0611# => '0' & O"331",
    8#0612# => '0' & O"704",
    8#0613# => '1' & O"264",
    8#0614# => '1' & O"007",
    8#0615# => '1' & O"364",
    8#0616# => '1' & O"137",
    8#0617# => '0' & O"424",
    8#0620# => '1' & O"117",
    8#0621# => '0' & O"146",
    8#0622# => '1' & O"637",
    8#0623# => '0' & O"250",
    8#0624# => '0' & O"612",
    8#0625# => '0' & O"114",
    8#0626# => '0' & O"416",
    8#0627# => '0' & O"074",
    8#0630# => '0' & O"454",
    8#0631# => '1' & O"133",
    8#0632# => '1' & O"662",
    8#0633# => '1' & O"414",
    8#0634# => '0' & O"642",
    8#0635# => '1' & O"177",
    8#0636# => '0' & O"546",
    8#0637# => '0' & O"250",
    8#0640# => '1' & O"637",
    8#0641# => '1' & O"324",
    8#0642# => '1' & O"507",
    8#0643# => '1' & O"273",
    8#0644# => '0' & O"014",
    8#0645# => '0' & O"542",
    8#0646# => '0' & O"542",
    8#0647# => '1' & O"247",
    8#0650# => '1' & O"020",
    8#0651# => '0' & O"542",
    8#0652# => '1' & O"263",
    8#0653# => '0' & O"420",
    8#0654# => '0' & O"542",
    8#0655# => '0' & O"567",
    8#0656# => '0' & O"620",
    8#0657# => '1' & O"656",
    8#0660# => '0' & O"250",
    8#0661# => '1' & O"652",
    8#0662# => '1' & O"044",
    8#0663# => '1' & O"557",
    8#0664# => '0' & O"424",
    8#0665# => '1' & O"117",
    8#0666# => '1' & O"613",
    8#0667# => '0' & O"621",
    8#0670# => '1' & O"701",
    8#0671# => '0' & O"250",
    8#0672# => '1' & O"264",
    8#0673# => '0' & O"420",
    8#0674# => '0' & O"542",
    8#0675# => '0' & O"157",
    8#0676# => '1' & O"661",
    8#0677# => '0' & O"224",
    8#0700# => '1' & O"713",
    8#0701# => '0' & O"061",
    8#0702# => '0' & O"214",
    8#0703# => '0' & O"230",
    8#0704# => '0' & O"132",
    8#0705# => '1' & O"707",
    8#0706# => '1' & O"732",
    8#0707# => '0' & O"061",
    8#0710# => '0' & O"347",
    8#0711# => '1' & O"024",
    8#0712# => '0' & O"137",
    8#0713# => '0' & O"324",
    8#0714# => '1' & O"243",
    8#0715# => '1' & O"207",
    8#0716# => '0' & O"030",
    8#0717# => '0' & O"564",
    8#0720# => '0' & O"663",
    8#0721# => '0' & O"164",
    8#0722# => '1' & O"543",
    8#0723# => '1' & O"044",
    8#0724# => '0' & O"620",
    8#0725# => '1' & O"656",
    8#0726# => '0' & O"250",
    8#0727# => '0' & O"422",
    8#0730# => '0' & O"014",
    8#0731# => '0' & O"602",
    8#0732# => '1' & O"656",
    8#0733# => '0' & O"250",
    8#0734# => '1' & O"656",
    8#0735# => '0' & O"621",
    8#0736# => '0' & O"461",
    8#0737# => '1' & O"025",
    8#0740# => '0' & O"624",
    8#0741# => '1' & O"323",
    8#0742# => '1' & O"065",
    8#0743# => '0' & O"624",
    8#0744# => '1' & O"077",
    8#0745# => '0' & O"676",
    8#0746# => '1' & O"117",
    8#0747# => '1' & O"025",
    8#0750# => '1' & O"656",
    8#0751# => '1' & O"735",
    8#0752# => '0' & O"564",
    8#0753# => '0' & O"117",
    8#0754# => '1' & O"044",
    8#0755# => '0' & O"620",
    8#0756# => '0' & O"000",
    8#0757# => '0' & O"336",
    8#0760# => '0' & O"620",
    8#0761# => '0' & O"061",
    8#0762# => '1' & O"701",
    8#0763# => '1' & O"124",
    8#0764# => '0' & O"533",
    8#0765# => '0' & O"704",
    8#0766# => '0' & O"347",
    8#0767# => '0' & O"564",
    8#0770# => '0' & O"643",
    8#0771# => '0' & O"250",
    8#0772# => '0' & O"624",
    8#0773# => '0' & O"013",
    8#0774# => '0' & O"332",
    8#0775# => '0' & O"772",
    8#0776# => '0' & O"250",
    8#0777# => '1' & O"701",
    8#1000# => '0' & O"321",
    8#1001# => '1' & O"767",
    8#1002# => '0' & O"646",
    8#1003# => '0' & O"447",
    8#1004# => '0' & O"176",
    8#1005# => '0' & O"447",
    8#1006# => '1' & O"124",
    8#1007# => '0' & O"353",
    8#1010# => '0' & O"204",
    8#1011# => '0' & O"616",
    8#1012# => '1' & O"224",
    8#1013# => '0' & O"363",
    8#1014# => '1' & O"356",
    8#1015# => '1' & O"506",
    8#1016# => '1' & O"316",
    8#1017# => '0' & O"576",
    8#1020# => '1' & O"620",
    8#1021# => '1' & O"364",
    8#1022# => '1' & O"143",
    8#1023# => '1' & O"261",
    8#1024# => '1' & O"701",
    8#1025# => '1' & O"056",
    8#1026# => '0' & O"343",
    8#1027# => '0' & O"450",
    8#1030# => '1' & O"656",
    8#1031# => '1' & O"204",
    8#1032# => '1' & O"414",
    8#1033# => '0' & O"043",
    8#1034# => '1' & O"220",
    8#1035# => '0' & O"621",
    8#1036# => '1' & O"521",
    8#1037# => '0' & O"650",
    8#1040# => '0' & O"450",
    8#1041# => '1' & O"656",
    8#1042# => '1' & O"037",
    8#1043# => '1' & O"264",
    8#1044# => '1' & O"343",
    8#1045# => '0' & O"621",
    8#1046# => '0' & O"565",
    8#1047# => '1' & O"521",
    8#1050# => '0' & O"650",
    8#1051# => '1' & O"176",
    8#1052# => '0' & O"467",
    8#1053# => '1' & O"146",
    8#1054# => '0' & O"137",
    8#1055# => '0' & O"013",
    8#1056# => '0' & O"316",
    8#1057# => '1' & O"414",
    8#1060# => '0' & O"430",
    8#1061# => '0' & O"752",
    8#1062# => '0' & O"060",
    8#1063# => '0' & O"167",
    8#1064# => '1' & O"364",
    8#1065# => '0' & O"477",
    8#1066# => '0' & O"250",
    8#1067# => '0' & O"064",
    8#1070# => '0' & O"220",
    8#1071# => '0' & O"000",
    8#1072# => '1' & O"656",
    8#1073# => '1' & O"037",
    8#1074# => '0' & O"524",
    8#1075# => '0' & O"407",
    8#1076# => '1' & O"764",
    8#1077# => '0' & O"047",
    8#1100# => '0' & O"000",
    8#1101# => '1' & O"620",
    8#1102# => '0' & O"216",
    8#1103# => '0' & O"376",
    8#1104# => '0' & O"115",
    8#1105# => '1' & O"701",
    8#1106# => '0' & O"404",
    8#1107# => '0' & O"343",
    8#1110# => '0' & O"000",
    8#1111# => '1' & O"124",
    8#1112# => '0' & O"467",
    8#1113# => '1' & O"144",
    8#1114# => '0' & O"503",
    8#1115# => '1' & O"656",
    8#1116# => '0' & O"450",
    8#1117# => '1' & O"656",
    8#1120# => '0' & O"764",
    8#1121# => '1' & O"413",
    8#1122# => '1' & O"521",
    8#1123# => '1' & O"701",
    8#1124# => '1' & O"124",
    8#1125# => '0' & O"413",
    8#1126# => '1' & O"656",
    8#1127# => '1' & O"224",
    8#1130# => '1' & O"003",
    8#1131# => '0' & O"372",
    8#1132# => '0' & O"616",
    8#1133# => '1' & O"364",
    8#1134# => '0' & O"653",
    8#1135# => '0' & O"144",
    8#1136# => '0' & O"244",
    8#1137# => '1' & O"103",
    8#1140# => '1' & O"261",
    8#1141# => '1' & O"015",
    8#1142# => '0' & O"014",
    8#1143# => '1' & O"527",
    8#1144# => '1' & O"220",
    8#1145# => '0' & O"164",
    8#1146# => '0' & O"257",
    8#1147# => '0' & O"000",
    8#1150# => '0' & O"104",
    8#1151# => '1' & O"077",
    8#1152# => '1' & O"364",
    8#1153# => '0' & O"107",
    8#1154# => '0' & O"416",
    8#1155# => '0' & O"034",
    8#1156# => '0' & O"054",
    8#1157# => '0' & O"663",
    8#1160# => '0' & O"714",
    8#1161# => '1' & O"642",
    8#1162# => '0' & O"250",
    8#1163# => '1' & O"656",
    8#1164# => '1' & O"261",
    8#1165# => '0' & O"621",
    8#1166# => '0' & O"117",
    8#1167# => '0' & O"000",
    8#1170# => '0' & O"000",
    8#1171# => '1' & O"364",
    8#1172# => '1' & O"137",
    8#1173# => '0' & O"104",
    8#1174# => '0' & O"573",
    8#1175# => '1' & O"656",
    8#1176# => '0' & O"164",
    8#1177# => '0' & O"237",
    8#1200# => '0' & O"376",
    8#1201# => '0' & O"616",
    8#1202# => '0' & O"343",
    8#1203# => '0' & O"250",
    8#1204# => '1' & O"656",
    8#1205# => '0' & O"250",
    8#1206# => '1' & O"443",
    8#1207# => '0' & O"220",
    8#1210# => '0' & O"424",
    8#1211# => '1' & O"063",
    8#1212# => '0' & O"321",
    8#1213# => '1' & O"037",
    8#1214# => '0' & O"161",
    8#1215# => '1' & O"037",
    8#1216# => '0' & O"144",
    8#1217# => '0' & O"204",
    8#1220# => '1' & O"056",
    8#1221# => '0' & O"316",
    8#1222# => '0' & O"752",
    8#1223# => '1' & O"414",
    8#1224# => '0' & O"230",
    8#1225# => '0' & O"124",
    8#1226# => '1' & O"143",
    8#1227# => '0' & O"130",
    8#1230# => '1' & O"160",
    8#1231# => '0' & O"224",
    8#1232# => '1' & O"447",
    8#1233# => '1' & O"370",
    8#1234# => '0' & O"124",
    8#1235# => '1' & O"443",
    8#1236# => '1' & O"656",
    8#1237# => '0' & O"650",
    8#1240# => '1' & O"656",
    8#1241# => '1' & O"370",
    8#1242# => '0' & O"450",
    8#1243# => '0' & O"216",
    8#1244# => '1' & O"443",
    8#1245# => '0' & O"161",
    8#1246# => '0' & O"450",
    8#1247# => '0' & O"572",
    8#1250# => '0' & O"672",
    8#1251# => '1' & O"367",
    8#1252# => '1' & O"307",
    8#1253# => '0' & O"000",
    8#1254# => '0' & O"304",
    8#1255# => '1' & O"344",
    8#1256# => '1' & O"044",
    8#1257# => '0' & O"060",
    8#1260# => '0' & O"000",
    8#1261# => '0' & O"372",
    8#1262# => '0' & O"672",
    8#1263# => '1' & O"343",
    8#1264# => '0' & O"572",
    8#1265# => '0' & O"172",
    8#1266# => '1' & O"347",
    8#1267# => '0' & O"572",
    8#1270# => '0' & O"321",
    8#1271# => '0' & O"316",
    8#1272# => '0' & O"742",
    8#1273# => '0' & O"105",
    8#1274# => '0' & O"625",
    8#1275# => '1' & O"376",
    8#1276# => '1' & O"071",
    8#1277# => '0' & O"321",
    8#1300# => '0' & O"650",
    8#1301# => '0' & O"450",
    8#1302# => '1' & O"656",
    8#1303# => '0' & O"651",
    8#1304# => '0' & O"164",
    8#1305# => '1' & O"007",
    8#1306# => '0' & O"216",
    8#1307# => '1' & O"360",
    8#1310# => '0' & O"220",
    8#1311# => '0' & O"124",
    8#1312# => '1' & O"433",
    8#1313# => '0' & O"216",
    8#1314# => '0' & O"456",
    8#1315# => '0' & O"650",
    8#1316# => '1' & O"656",
    8#1317# => '1' & O"360",
    8#1320# => '0' & O"450",
    8#1321# => '1' & O"456",
    8#1322# => '1' & O"217",
    8#1323# => '0' & O"000",
    8#1324# => '0' & O"620",
    8#1325# => '0' & O"602",
    8#1326# => '1' & O"015",
    8#1327# => '0' & O"621",
    8#1330# => '0' & O"565",
    8#1331# => '1' & O"056",
    8#1332# => '1' & O"250",
    8#1333# => '1' & O"356",
    8#1334# => '0' & O"014",
    8#1335# => '0' & O"602",
    8#1336# => '0' & O"316",
    8#1337# => '1' & O"552",
    8#1340# => '0' & O"217",
    8#1341# => '0' & O"216",
    8#1342# => '0' & O"755",
    8#1343# => '0' & O"650",
    8#1344# => '1' & O"204",
    8#1345# => '0' & O"424",
    8#1346# => '0' & O"767",
    8#1347# => '0' & O"156",
    8#1350# => '1' & O"227",
    8#1351# => '1' & O"156",
    8#1352# => '1' & O"667",
    8#1353# => '0' & O"450",
    8#1354# => '1' & O"037",
    8#1355# => '0' & O"456",
    8#1356# => '0' & O"764",
    8#1357# => '1' & O"043",
    8#1360# => '0' & O"620",
    8#1361# => '1' & O"456",
    8#1362# => '0' & O"524",
    8#1363# => '1' & O"043",
    8#1364# => '0' & O"271",
    8#1365# => '0' & O"105",
    8#1366# => '0' & O"316",
    8#1367# => '1' & O"414",
    8#1370# => '0' & O"130",
    8#1371# => '1' & O"030",
    8#1372# => '0' & O"424",
    8#1373# => '0' & O"003",
    8#1374# => '0' & O"161",
    8#1375# => '0' & O"271",
    8#1376# => '0' & O"745",
    8#1377# => '1' & O"037",
    8#1400# => '1' & O"767",
    8#1401# => '1' & O"656",
    8#1402# => '1' & O"414",
    8#1403# => '0' & O"130",
    8#1404# => '0' & O"752",
    8#1405# => '1' & O"160",
    8#1406# => '0' & O"250",
    8#1407# => '1' & O"656",
    8#1410# => '0' & O"250",
    8#1411# => '0' & O"621",
    8#1412# => '0' & O"250",
    8#1413# => '0' & O"572",
    8#1414# => '1' & O"017",
    8#1415# => '0' & O"250",
    8#1416# => '1' & O"360",
    8#1417# => '1' & O"037",
    8#1420# => '1' & O"275",
    8#1421# => '0' & O"621",
    8#1422# => '1' & O"264",
    8#1423# => '0' & O"377",
    8#1424# => '0' & O"621",
    8#1425# => '1' & O"525",
    8#1426# => '1' & O"450",
    8#1427# => '1' & O"037",
    8#1430# => '1' & O"705",
    8#1431# => '1' & O"124",
    8#1432# => '1' & O"237",
    8#1433# => '1' & O"056",
    8#1434# => '1' & O"146",
    8#1435# => '0' & O"327",
    8#1436# => '1' & O"414",
    8#1437# => '1' & O"356",
    8#1440# => '0' & O"316",
    8#1441# => '1' & O"742",
    8#1442# => '0' & O"562",
    8#1443# => '0' & O"230",
    8#1444# => '0' & O"327",
    8#1445# => '0' & O"747",
    8#1446# => '0' & O"542",
    8#1447# => '0' & O"742",
    8#1450# => '1' & O"447",
    8#1451# => '0' & O"250",
    8#1452# => '1' & O"545",
    8#1453# => '1' & O"515",
    8#1454# => '0' & O"305",
    8#1455# => '0' & O"275",
    8#1456# => '1' & O"453",
    8#1457# => '1' & O"364",
    8#1460# => '0' & O"167",
    8#1461# => '0' & O"164",
    8#1462# => '1' & O"453",
    8#1463# => '0' & O"123",
    8#1464# => '0' & O"000",
    8#1465# => '0' & O"312",
    8#1466# => '1' & O"204",
    8#1467# => '1' & O"056",
    8#1470# => '0' & O"220",
    8#1471# => '0' & O"572",
    8#1472# => '0' & O"373",
    8#1473# => '1' & O"601",
    8#1474# => '1' & O"515",
    8#1475# => '0' & O"647",
    8#1476# => '0' & O"250",
    8#1477# => '0' & O"656",
    8#1500# => '1' & O"413",
    8#1501# => '1' & O"605",
    8#1502# => '0' & O"275",
    8#1503# => '0' & O"647",
    8#1504# => '0' & O"000",
    8#1505# => '1' & O"633",
    8#1506# => '1' & O"356",
    8#1507# => '0' & O"014",
    8#1510# => '0' & O"602",
    8#1511# => '0' & O"416",
    8#1512# => '0' & O"074",
    8#1513# => '1' & O"454",
    8#1514# => '0' & O"447",
    8#1515# => '1' & O"656",
    8#1516# => '1' & O"160",
    8#1517# => '1' & O"656",
    8#1520# => '0' & O"060",
    8#1521# => '0' & O"000",
    8#1522# => '0' & O"624",
    8#1523# => '0' & O"143",
    8#1524# => '0' & O"621",
    8#1525# => '0' & O"561",
    8#1526# => '1' & O"264",
    8#1527# => '0' & O"420",
    8#1530# => '1' & O"364",
    8#1531# => '1' & O"143",
    8#1532# => '0' & O"564",
    8#1533# => '0' & O"643",
    8#1534# => '0' & O"420",
    8#1535# => '0' & O"124",
    8#1536# => '0' & O"603",
    8#1537# => '1' & O"144",
    8#1540# => '0' & O"224",
    8#1541# => '1' & O"267",
    8#1542# => '1' & O"037",
    8#1543# => '0' & O"000",
    8#1544# => '1' & O"220",
    8#1545# => '0' & O"572",
    8#1546# => '1' & O"337",
    8#1547# => '1' & O"601",
    8#1550# => '0' & O"541",
    8#1551# => '1' & O"361",
    8#1552# => '1' & O"370",
    8#1553# => '1' & O"656",
    8#1554# => '1' & O"360",
    8#1555# => '1' & O"656",
    8#1556# => '1' & O"037",
    8#1557# => '0' & O"564",
    8#1560# => '1' & O"073",
    8#1561# => '0' & O"572",
    8#1562# => '0' & O"627",
    8#1563# => '0' & O"431",
    8#1564# => '0' & O"250",
    8#1565# => '0' & O"724",
    8#1566# => '1' & O"033",
    8#1567# => '0' & O"450",
    8#1570# => '1' & O"033",
    8#1571# => '0' & O"621",
    8#1572# => '0' & O"561",
    8#1573# => '1' & O"525",
    8#1574# => '0' & O"656",
    8#1575# => '1' & O"413",
    8#1576# => '1' & O"356",
    8#1577# => '1' & O"414",
    8#1600# => '1' & O"742",
    8#1601# => '0' & O"275",
    8#1602# => '1' & O"037",
    8#1603# => '0' & O"572",
    8#1604# => '1' & O"317",
    8#1605# => '0' & O"723",
    8#1606# => '1' & O"370",
    8#1607# => '0' & O"220",
    8#1610# => '1' & O"275",
    8#1611# => '0' & O"305",
    8#1612# => '0' & O"036",
    8#1613# => '1' & O"067",
    8#1614# => '0' & O"576",
    8#1615# => '1' & O"275",
    8#1616# => '0' & O"450",
    8#1617# => '0' & O"616",
    8#1620# => '0' & O"551",
    8#1621# => '1' & O"224",
    8#1622# => '1' & O"163",
    8#1623# => '0' & O"675",
    8#1624# => '0' & O"676",
    8#1625# => '1' & O"163",
    8#1626# => '0' & O"305",
    8#1627# => '1' & O"256",
    8#1630# => '1' & O"176",
    8#1631# => '1' & O"157",
    8#1632# => '0' & O"576",
    8#1633# => '0' & O"541",
    8#1634# => '1' & O"656",
    8#1635# => '0' & O"616",
    8#1636# => '0' & O"250",
    8#1637# => '0' & O"614",
    8#1640# => '0' & O"742",
    8#1641# => '0' & O"542",
    8#1642# => '0' & O"233",
    8#1643# => '0' & O"250",
    8#1644# => '1' & O"752",
    8#1645# => '1' & O"752",
    8#1646# => '0' & O"261",
    8#1647# => '0' & O"724",
    8#1650# => '1' & O"257",
    8#1651# => '1' & O"056",
    8#1652# => '0' & O"450",
    8#1653# => '1' & O"104",
    8#1654# => '0' & O"173",
    8#1655# => '0' & O"364",
    8#1656# => '1' & O"447",
    8#1657# => '0' & O"304",
    8#1660# => '1' & O"304",
    8#1661# => '1' & O"004",
    8#1662# => '0' & O"060",
    8#1663# => '0' & O"572",
    8#1664# => '0' & O"707",
    8#1665# => '0' & O"431",
    8#1666# => '0' & O"067",
    8#1667# => '0' & O"572",
    8#1670# => '0' & O"347",
    8#1671# => '1' & O"601",
    8#1672# => '1' & O"571",
    8#1673# => '0' & O"647",
    8#1674# => '1' & O"364",
    8#1675# => '0' & O"107",
    8#1676# => '0' & O"000",
    8#1677# => '1' & O"275",
    8#1700# => '0' & O"551",
    8#1701# => '0' & O"675",
    8#1702# => '0' & O"250",
    8#1703# => '1' & O"414",
    8#1704# => '0' & O"302",
    8#1705# => '0' & O"250",
    8#1706# => '0' & O"064",
    8#1707# => '0' & O"504",
    8#1710# => '0' & O"337",
    8#1711# => '0' & O"250",
    8#1712# => '1' & O"361",
    8#1713# => '1' & O"144",
    8#1714# => '1' & O"224",
    8#1715# => '1' & O"037",
    8#1716# => '0' & O"650",
    8#1717# => '0' & O"450",
    8#1720# => '1' & O"376",
    8#1721# => '1' & O"656",
    8#1722# => '1' & O"037",
    8#1723# => '1' & O"364",
    8#1724# => '0' & O"477",
    8#1725# => '0' & O"424",
    8#1726# => '1' & O"673",
    8#1727# => '0' & O"020",
    8#1730# => '0' & O"000",
    8#1731# => '0' & O"164",
    8#1732# => '0' & O"463",
    8#1733# => '0' & O"224",
    8#1734# => '0' & O"567",
    8#1735# => '0' & O"577",
    8#1736# => '1' & O"364",
    8#1737# => '1' & O"137",
    8#1740# => '0' & O"250",
    8#1741# => '0' & O"616",
    8#1742# => '1' & O"370",
    8#1743# => '1' & O"656",
    8#1744# => '1' & O"360",
    8#1745# => '0' & O"060",
    8#1746# => '1' & O"525",
    8#1747# => '1' & O"705",
    8#1750# => '0' & O"250",
    8#1751# => '0' & O"332",
    8#1752# => '0' & O"204",
    8#1753# => '0' & O"250",
    8#1754# => '0' & O"343",
    8#1755# => '0' & O"000",
    8#1756# => '0' & O"624",
    8#1757# => '1' & O"267",
    8#1760# => '1' & O"537",
    8#1761# => '0' & O"644",
    8#1762# => '0' & O"244",
    8#1763# => '0' & O"444",
    8#1764# => '0' & O"144",
    8#1765# => '1' & O"267",
    8#1766# => '1' & O"275",
    8#1767# => '0' & O"250",
    8#1770# => '1' & O"656",
    8#1771# => '0' & O"250",
    8#1772# => '0' & O"014",
    8#1773# => '0' & O"602",
    8#1774# => '1' & O"656",
    8#1775# => '0' & O"416",
    8#1776# => '0' & O"074",
    8#1777# => '1' & O"354",
    8#2000# => '0' & O"060",
    8#2001# => '1' & O"151",
    8#2002# => '0' & O"471",
    8#2003# => '0' & O"650",
    8#2004# => '1' & O"135",
    8#2005# => '0' & O"450",
    8#2006# => '0' & O"305",
    8#2007# => '1' & O"341",
    8#2010# => '0' & O"616",
    8#2011# => '0' & O"471",
    8#2012# => '1' & O"345",
    8#2013# => '0' & O"575",
    8#2014# => '0' & O"415",
    8#2015# => '1' & O"335",
    8#2016# => '1' & O"131",
    8#2017# => '0' & O"624",
    8#2020# => '1' & O"233",
    8#2021# => '0' & O"605",
    8#2022# => '0' & O"475",
    8#2023# => '0' & O"565",
    8#2024# => '0' & O"305",
    8#2025# => '1' & O"321",
    8#2026# => '0' & O"616",
    8#2027# => '1' & O"341",
    8#2030# => '0' & O"471",
    8#2031# => '0' & O"475",
    8#2032# => '0' & O"305",
    8#2033# => '1' & O"331",
    8#2034# => '0' & O"616",
    8#2035# => '1' & O"335",
    8#2036# => '0' & O"471",
    8#2037# => '0' & O"650",
    8#2040# => '1' & O"131",
    8#2041# => '1' & O"345",
    8#2042# => '0' & O"415",
    8#2043# => '0' & O"450",
    8#2044# => '1' & O"043",
    8#2045# => '1' & O"364",
    8#2046# => '0' & O"263",
    8#2047# => '0' & O"724",
    8#2050# => '1' & O"443",
    8#2051# => '0' & O"572",
    8#2052# => '0' & O"172",
    8#2053# => '1' & O"443",
    8#2054# => '1' & O"215",
    8#2055# => '1' & O"331",
    8#2056# => '0' & O"475",
    8#2057# => '1' & O"215",
    8#2060# => '1' & O"033",
    8#2061# => '1' & O"656",
    8#2062# => '1' & O"217",
    8#2063# => '0' & O"621",
    8#2064# => '0' & O"444",
    8#2065# => '0' & O"704",
    8#2066# => '0' & O"561",
    8#2067# => '0' & O"565",
    8#2070# => '0' & O"033",
    8#2071# => '0' & O"424",
    8#2072# => '0' & O"453",
    8#2073# => '0' & O"444",
    8#2074# => '1' & O"215",
    8#2075# => '1' & O"345",
    8#2076# => '1' & O"356",
    8#2077# => '1' & O"742",
    8#2100# => '1' & O"507",
    8#2101# => '1' & O"364",
    8#2102# => '0' & O"107",
    8#2103# => '1' & O"364",
    8#2104# => '0' & O"167",
    8#2105# => '1' & O"161",
    8#2106# => '0' & O"604",
    8#2107# => '1' & O"313",
    8#2110# => '0' & O"764",
    8#2111# => '1' & O"527",
    8#2112# => '0' & O"450",
    8#2113# => '1' & O"141",
    8#2114# => '1' & O"303",
    8#2115# => '0' & O"237",
    8#2116# => '1' & O"220",
    8#2117# => '0' & O"650",
    8#2120# => '0' & O"450",
    8#2121# => '0' & O"060",
    8#2122# => '1' & O"267",
    8#2123# => '1' & O"201",
    8#2124# => '1' & O"331",
    8#2125# => '0' & O"704",
    8#2126# => '1' & O"507",
    8#2127# => '1' & O"151",
    8#2130# => '1' & O"215",
    8#2131# => '1' & O"341",
    8#2132# => '0' & O"404",
    8#2133# => '1' & O"507",
    8#2134# => '0' & O"420",
    8#2135# => '0' & O"564",
    8#2136# => '0' & O"757",
    8#2137# => '0' & O"176",
    8#2140# => '1' & O"373",
    8#2141# => '0' & O"646",
    8#2142# => '1' & O"373",
    8#2143# => '0' & O"060",
    8#2144# => '1' & O"220",
    8#2145# => '1' & O"356",
    8#2146# => '1' & O"742",
    8#2147# => '1' & O"131",
    8#2150# => '1' & O"771",
    8#2151# => '0' & O"475",
    8#2152# => '0' & O"565",
    8#2153# => '0' & O"305",
    8#2154# => '1' & O"331",
    8#2155# => '0' & O"616",
    8#2156# => '0' & O"471",
    8#2157# => '1' & O"345",
    8#2160# => '0' & O"415",
    8#2161# => '1' & O"325",
    8#2162# => '1' & O"131",
    8#2163# => '0' & O"475",
    8#2164# => '0' & O"033",
    8#2165# => '1' & O"341",
    8#2166# => '0' & O"475",
    8#2167# => '1' & O"141",
    8#2170# => '0' & O"456",
    8#2171# => '0' & O"475",
    8#2172# => '0' & O"216",
    8#2173# => '1' & O"656",
    8#2174# => '0' & O"415",
    8#2175# => '0' & O"424",
    8#2176# => '1' & O"007",
    8#2177# => '0' & O"336",
    8#2200# => '1' & O"171",
    8#2201# => '0' & O"405",
    8#2202# => '0' & O"724",
    8#2203# => '1' & O"037",
    8#2204# => '0' & O"744",
    8#2205# => '0' & O"733",
    8#2206# => '1' & O"341",
    8#2207# => '0' & O"220",
    8#2210# => '0' & O"305",
    8#2211# => '1' & O"341",
    8#2212# => '0' & O"616",
    8#2213# => '1' & O"331",
    8#2214# => '0' & O"471",
    8#2215# => '1' & O"345",
    8#2216# => '0' & O"415",
    8#2217# => '1' & O"321",
    8#2220# => '1' & O"131",
    8#2221# => '0' & O"724",
    8#2222# => '0' & O"007",
    8#2223# => '0' & O"475",
    8#2224# => '1' & O"656",
    8#2225# => '0' & O"733",
    8#2226# => '0' & O"376",
    8#2227# => '1' & O"220",
    8#2230# => '0' & O"564",
    8#2231# => '0' & O"643",
    8#2232# => '0' & O"564",
    8#2233# => '1' & O"073",
    8#2234# => '0' & O"764",
    8#2235# => '1' & O"707",
    8#2236# => '0' & O"164",
    8#2237# => '0' & O"257",
    8#2240# => '0' & O"650",
    8#2241# => '1' & O"656",
    8#2242# => '0' & O"450",
    8#2243# => '0' & O"616",
    8#2244# => '1' & O"414",
    8#2245# => '0' & O"060",
    8#2246# => '0' & O"424",
    8#2247# => '1' & O"617",
    8#2250# => '0' & O"733",
    8#2251# => '0' & O"344",
    8#2252# => '1' & O"344",
    8#2253# => '1' & O"004",
    8#2254# => '0' & O"060",
    8#2255# => '0' & O"621",
    8#2256# => '0' & O"441",
    8#2257# => '0' & O"450",
    8#2260# => '1' & O"056",
    8#2261# => '0' & O"064",
    8#2262# => '0' & O"364",
    8#2263# => '0' & O"347",
    8#2264# => '0' & O"542",
    8#2265# => '0' & O"542",
    8#2266# => '0' & O"542",
    8#2267# => '0' & O"542",
    8#2270# => '0' & O"542",
    8#2271# => '0' & O"516",
    8#2272# => '1' & O"160",
    8#2273# => '0' & O"000",
    8#2274# => '1' & O"370",
    8#2275# => '0' & O"060",
    8#2276# => '0' & O"620",
    8#2277# => '0' & O"724",
    8#2300# => '0' & O"347",
    8#2301# => '0' & O"744",
    8#2302# => '1' & O"151",
    8#2303# => '1' & O"215",
    8#2304# => '1' & O"321",
    8#2305# => '1' & O"656",
    8#2306# => '0' & O"650",
    8#2307# => '1' & O"477",
    8#2310# => '0' & O"565",
    8#2311# => '0' & O"744",
    8#2312# => '1' & O"204",
    8#2313# => '1' & O"201",
    8#2314# => '1' & O"325",
    8#2315# => '1' & O"656",
    8#2316# => '0' & O"616",
    8#2317# => '0' & O"471",
    8#2320# => '1' & O"370",
    8#2321# => '1' & O"656",
    8#2322# => '0' & O"624",
    8#2323# => '1' & O"527",
    8#2324# => '0' & O"376",
    8#2325# => '1' & O"135",
    8#2326# => '0' & O"405",
    8#2327# => '1' & O"360",
    8#2330# => '1' & O"224",
    8#2331# => '1' & O"377",
    8#2332# => '0' & O"724",
    8#2333# => '0' & O"517",
    8#2334# => '0' & O"424",
    8#2335# => '0' & O"537",
    8#2336# => '1' & O"151",
    8#2337# => '1' & O"215",
    8#2340# => '1' & O"335",
    8#2341# => '1' & O"244",
    8#2342# => '1' & O"467",
    8#2343# => '0' & O"605",
    8#2344# => '0' & O"724",
    8#2345# => '1' & O"747",
    8#2346# => '0' & O"744",
    8#2347# => '0' & O"123",
    8#2350# => '1' & O"245",
    8#2351# => '0' & O"621",
    8#2352# => '0' & O"561",
    8#2353# => '0' & O"565",
    8#2354# => '0' & O"704",
    8#2355# => '0' & O"305",
    8#2356# => '1' & O"345",
    8#2357# => '0' & O"624",
    8#2360# => '0' & O"627",
    8#2361# => '0' & O"575",
    8#2362# => '0' & O"475",
    8#2363# => '0' & O"565",
    8#2364# => '0' & O"305",
    8#2365# => '1' & O"331",
    8#2366# => '0' & O"475",
    8#2367# => '0' & O"305",
    8#2370# => '0' & O"727",
    8#2371# => '0' & O"650",
    8#2372# => '0' & O"415",
    8#2373# => '0' & O"450",
    8#2374# => '1' & O"141",
    8#2375# => '1' & O"037",
    8#2376# => '0' & O"676",
    8#2377# => '1' & O"373",
    8#2400# => '0' & O"556",
    8#2401# => '0' & O"354",
    8#2402# => '0' & O"023",
    8#2403# => '0' & O"043",
    8#2404# => '0' & O"724",
    8#2405# => '0' & O"037",
    8#2406# => '0' & O"034",
    8#2407# => '1' & O"122",
    8#2410# => '1' & O"352",
    8#2411# => '1' & O"056",
    8#2412# => '0' & O"553",
    8#2413# => '0' & O"322",
    8#2414# => '0' & O"562",
    8#2415# => '0' & O"332",
    8#2416# => '1' & O"612",
    8#2417# => '1' & O"513",
    8#2420# => '0' & O"316",
    8#2421# => '0' & O"616",
    8#2422# => '1' & O"414",
    8#2423# => '0' & O"452",
    8#2424# => '0' & O"612",
    8#2425# => '0' & O"672",
    8#2426# => '0' & O"153",
    8#2427# => '0' & O"252",
    8#2430# => '0' & O"572",
    8#2431# => '0' & O"057",
    8#2432# => '1' & O"652",
    8#2433# => '0' & O"616",
    8#2434# => '1' & O"443",
    8#2435# => '1' & O"414",
    8#2436# => '0' & O"056",
    8#2437# => '0' & O"144",
    8#2440# => '0' & O"244",
    8#2441# => '1' & O"564",
    8#2442# => '1' & O"233",
    8#2443# => '1' & O"256",
    8#2444# => '1' & O"443",
    8#2445# => '1' & O"025",
    8#2446# => '0' & O"224",
    8#2447# => '0' & O"757",
    8#2450# => '0' & O"172",
    8#2451# => '0' & O"757",
    8#2452# => '0' & O"730",
    8#2453# => '0' & O"547",
    8#2454# => '1' & O"471",
    8#2455# => '0' & O"625",
    8#2456# => '0' & O"744",
    8#2457# => '0' & O"224",
    8#2460# => '0' & O"447",
    8#2461# => '0' & O"704",
    8#2462# => '0' & O"447",
    8#2463# => '1' & O"025",
    8#2464# => '0' & O"224",
    8#2465# => '0' & O"367",
    8#2466# => '0' & O"172",
    8#2467# => '0' & O"367",
    8#2470# => '0' & O"630",
    8#2471# => '0' & O"547",
    8#2472# => '1' & O"004",
    8#2473# => '1' & O"264",
    8#2474# => '0' & O"220",
    8#2475# => '0' & O"250",
    8#2476# => '0' & O"625",
    8#2477# => '1' & O"015",
    8#2500# => '0' & O"561",
    8#2501# => '0' & O"650",
    8#2502# => '0' & O"475",
    8#2503# => '1' & O"013",
    8#2504# => '0' & O"000",
    8#2505# => '1' & O"025",
    8#2506# => '1' & O"317",
    8#2507# => '0' & O"602",
    8#2510# => '0' & O"653",
    8#2511# => '0' & O"444",
    8#2512# => '0' & O"561",
    8#2513# => '1' & O"250",
    8#2514# => '0' & O"465",
    8#2515# => '1' & O"164",
    8#2516# => '1' & O"247",
    8#2517# => '0' & O"252",
    8#2520# => '0' & O"314",
    8#2521# => '0' & O"173",
    8#2522# => '1' & O"025",
    8#2523# => '1' & O"053",
    8#2524# => '0' & O"000",
    8#2525# => '0' & O"622",
    8#2526# => '1' & O"056",
    8#2527# => '1' & O"733",
    8#2530# => '0' & O"430",
    8#2531# => '0' & O"250",
    8#2532# => '0' & O"364",
    8#2533# => '0' & O"347",
    8#2534# => '0' & O"420",
    8#2535# => '0' & O"114",
    8#2536# => '1' & O"124",
    8#2537# => '1' & O"653",
    8#2540# => '1' & O"224",
    8#2541# => '0' & O"527",
    8#2542# => '0' & O"422",
    8#2543# => '0' & O"014",
    8#2544# => '0' & O"437",
    8#2545# => '1' & O"124",
    8#2546# => '1' & O"423",
    8#2547# => '0' & O"704",
    8#2550# => '1' & O"144",
    8#2551# => '1' & O"244",
    8#2552# => '1' & O"656",
    8#2553# => '0' & O"646",
    8#2554# => '0' & O"103",
    8#2555# => '0' & O"616",
    8#2556# => '0' & O"672",
    8#2557# => '0' & O"707",
    8#2560# => '1' & O"420",
    8#2561# => '0' & O"052",
    8#2562# => '1' & O"452",
    8#2563# => '1' & O"514",
    8#2564# => '0' & O"002",
    8#2565# => '1' & O"377",
    8#2566# => '1' & O"552",
    8#2567# => '0' & O"034",
    8#2570# => '0' & O"254",
    8#2571# => '1' & O"277",
    8#2572# => '1' & O"457",
    8#2573# => '0' & O"250",
    8#2574# => '0' & O"625",
    8#2575# => '0' & O"561",
    8#2576# => '0' & O"656",
    8#2577# => '1' & O"043",
    8#2600# => '0' & O"650",
    8#2601# => '0' & O"165",
    8#2602# => '1' & O"020",
    8#2603# => '0' & O"764",
    8#2604# => '1' & O"673",
    8#2605# => '0' & O"214",
    8#2606# => '0' & O"250",
    8#2607# => '0' & O"060",
    8#2610# => '0' & O"764",
    8#2611# => '1' & O"413",
    8#2612# => '0' & O"224",
    8#2613# => '1' & O"073",
    8#2614# => '0' & O"672",
    8#2615# => '1' & O"127",
    8#2616# => '0' & O"250",
    8#2617# => '0' & O"625",
    8#2620# => '1' & O"015",
    8#2621# => '0' & O"561",
    8#2622# => '0' & O"650",
    8#2623# => '1' & O"135",
    8#2624# => '1' & O"013",
    8#2625# => '0' & O"530",
    8#2626# => '0' & O"547",
    8#2627# => '0' & O"376",
    8#2630# => '0' & O"144",
    8#2631# => '0' & O"244",
    8#2632# => '1' & O"414",
    8#2633# => '0' & O"056",
    8#2634# => '1' & O"772",
    8#2635# => '1' & O"772",
    8#2636# => '0' & O"772",
    8#2637# => '0' & O"772",
    8#2640# => '0' & O"112",
    8#2641# => '1' & O"217",
    8#2642# => '1' & O"656",
    8#2643# => '1' & O"646",
    8#2644# => '0' & O"646",
    8#2645# => '1' & O"237",
    8#2646# => '1' & O"656",
    8#2647# => '1' & O"046",
    8#2650# => '0' & O"112",
    8#2651# => '1' & O"373",
    8#2652# => '1' & O"216",
    8#2653# => '1' & O"752",
    8#2654# => '0' & O"016",
    8#2655# => '1' & O"373",
    8#2656# => '1' & O"243",
    8#2657# => '0' & O"142",
    8#2660# => '1' & O"457",
    8#2661# => '0' & O"406",
    8#2662# => '0' & O"733",
    8#2663# => '0' & O"224",
    8#2664# => '1' & O"337",
    8#2665# => '0' & O"672",
    8#2666# => '0' & O"543",
    8#2667# => '0' & O"250",
    8#2670# => '0' & O"625",
    8#2671# => '1' & O"015",
    8#2672# => '0' & O"561",
    8#2673# => '0' & O"650",
    8#2674# => '1' & O"141",
    8#2675# => '1' & O"013",
    8#2676# => '1' & O"420",
    8#2677# => '0' & O"034",
    8#2700# => '0' & O"142",
    8#2701# => '1' & O"447",
    8#2702# => '0' & O"406",
    8#2703# => '0' & O"723",
    8#2704# => '1' & O"056",
    8#2705# => '0' & O"146",
    8#2706# => '1' & O"443",
    8#2707# => '0' & O"316",
    8#2710# => '0' & O"220",
    8#2711# => '0' & O"002",
    8#2712# => '1' & O"557",
    8#2713# => '1' & O"712",
    8#2714# => '1' & O"656",
    8#2715# => '1' & O"573",
    8#2716# => '0' & O"304",
    8#2717# => '1' & O"304",
    8#2720# => '1' & O"044",
    8#2721# => '0' & O"060",
    8#2722# => '0' & O"250",
    8#2723# => '0' & O"302",
    8#2724# => '0' & O"250",
    8#2725# => '0' & O"107",
    8#2726# => '0' & O"124",
    8#2727# => '0' & O"217",
    8#2730# => '1' & O"420",
    8#2731# => '1' & O"414",
    8#2732# => '1' & O"533",
    8#2733# => '1' & O"752",
    8#2734# => '0' & O"034",
    8#2735# => '1' & O"447",
    8#2736# => '1' & O"452",
    8#2737# => '0' & O"052",
    8#2740# => '1' & O"124",
    8#2741# => '0' & O"107",
    8#2742# => '0' & O"672",
    8#2743# => '0' & O"553",
    8#2744# => '0' & O"252",
    8#2745# => '0' & O"672",
    8#2746# => '0' & O"553",
    8#2747# => '1' & O"471",
    8#2750# => '0' & O"635",
    8#2751# => '1' & O"013",
    8#2752# => '1' & O"056",
    8#2753# => '1' & O"104",
    8#2754# => '0' & O"724",
    8#2755# => '1' & O"703",
    8#2756# => '0' & O"744",
    8#2757# => '0' & O"450",
    8#2760# => '1' & O"462",
    8#2761# => '1' & O"376",
    8#2762# => '0' & O"316",
    8#2763# => '0' & O"556",
    8#2764# => '0' & O"276",
    8#2765# => '0' & O"776",
    8#2766# => '0' & O"756",
    8#2767# => '0' & O"142",
    8#2770# => '0' & O"003",
    8#2771# => '0' & O"422",
    8#2772# => '0' & O"074",
    8#2773# => '1' & O"737",
    8#2774# => '1' & O"471",
    8#2775# => '0' & O"625",
    8#2776# => '1' & O"056",
    8#2777# => '0' & O"353",
    8#3000# => '1' & O"717",
    8#3001# => '1' & O"456",
    8#3002# => '0' & O"241",
    8#3003# => '0' & O"650",
    8#3004# => '0' & O"241",
    8#3005# => '0' & O"650",
    8#3006# => '1' & O"124",
    8#3007# => '0' & O"047",
    8#3010# => '1' & O"656",
    8#3011# => '0' & O"524",
    8#3012# => '0' & O"113",
    8#3013# => '0' & O"336",
    8#3014# => '1' & O"231",
    8#3015# => '0' & O"450",
    8#3016# => '1' & O"225",
    8#3017# => '1' & O"141",
    8#3020# => '0' & O"225",
    8#3021# => '0' & O"650",
    8#3022# => '1' & O"231",
    8#3023# => '0' & O"424",
    8#3024# => '0' & O"723",
    8#3025# => '1' & O"356",
    8#3026# => '1' & O"742",
    8#3027# => '0' & O"446",
    8#3030# => '1' & O"646",
    8#3031# => '0' & O"552",
    8#3032# => '1' & O"222",
    8#3033# => '0' & O"672",
    8#3034# => '0' & O"147",
    8#3035# => '1' & O"322",
    8#3036# => '0' & O"752",
    8#3037# => '0' & O"167",
    8#3040# => '1' & O"316",
    8#3041# => '1' & O"216",
    8#3042# => '0' & O"450",
    8#3043# => '1' & O"056",
    8#3044# => '0' & O"407",
    8#3045# => '1' & O"056",
    8#3046# => '0' & O"414",
    8#3047# => '1' & O"573",
    8#3050# => '0' & O"450",
    8#3051# => '1' & O"656",
    8#3052# => '0' & O"642",
    8#3053# => '0' & O"267",
    8#3054# => '0' & O"256",
    8#3055# => '0' & O"616",
    8#3056# => '0' & O"212",
    8#3057# => '1' & O"457",
    8#3060# => '0' & O"616",
    8#3061# => '0' & O"124",
    8#3062# => '0' & O"227",
    8#3063# => '0' & O"424",
    8#3064# => '0' & O"733",
    8#3065# => '0' & O"524",
    8#3066# => '0' & O"127",
    8#3067# => '0' & O"376",
    8#3070# => '1' & O"676",
    8#3071# => '0' & O"067",
    8#3072# => '1' & O"222",
    8#3073# => '1' & O"576",
    8#3074# => '0' & O"353",
    8#3075# => '0' & O"776",
    8#3076# => '1' & O"462",
    8#3077# => '0' & O"722",
    8#3100# => '1' & O"456",
    8#3101# => '0' & O"456",
    8#3102# => '1' & O"522",
    8#3103# => '0' & O"357",
    8#3104# => '0' & O"650",
    8#3105# => '1' & O"316",
    8#3106# => '1' & O"662",
    8#3107# => '1' & O"456",
    8#3110# => '0' & O"422",
    8#3111# => '0' & O"450",
    8#3112# => '1' & O"776",
    8#3113# => '1' & O"776",
    8#3114# => '0' & O"217",
    8#3115# => '0' & O"316",
    8#3116# => '0' & O"052",
    8#3117# => '1' & O"326",
    8#3120# => '1' & O"311",
    8#3121# => '0' & O"542",
    8#3122# => '0' & O"650",
    8#3123# => '1' & O"656",
    8#3124# => '0' & O"414",
    8#3125# => '1' & O"221",
    8#3126# => '0' & O"614",
    8#3127# => '1' & O"155",
    8#3130# => '1' & O"014",
    8#3131# => '1' & O"155",
    8#3132# => '0' & O"214",
    8#3133# => '1' & O"030",
    8#3134# => '1' & O"214",
    8#3135# => '1' & O"155",
    8#3136# => '1' & O"071",
    8#3137# => '1' & O"155",
    8#3140# => '1' & O"461",
    8#3141# => '0' & O"416",
    8#3142# => '1' & O"155",
    8#3143# => '0' & O"216",
    8#3144# => '1' & O"455",
    8#3145# => '1' & O"461",
    8#3146# => '1' & O"256",
    8#3147# => '1' & O"231",
    8#3150# => '1' & O"124",
    8#3151# => '0' & O"663",
    8#3152# => '0' & O"376",
    8#3153# => '1' & O"141",
    8#3154# => '1' & O"461",
    8#3155# => '1' & O"256",
    8#3156# => '1' & O"225",
    8#3157# => '0' & O"764",
    8#3160# => '1' & O"067",
    8#3161# => '0' & O"252",
    8#3162# => '1' & O"764",
    8#3163# => '0' & O"073",
    8#3164# => '0' & O"164",
    8#3165# => '1' & O"463",
    8#3166# => '1' & O"461",
    8#3167# => '1' & O"256",
    8#3170# => '1' & O"256",
    8#3171# => '1' & O"125",
    8#3172# => '1' & O"256",
    8#3173# => '1' & O"655",
    8#3174# => '1' & O"461",
    8#3175# => '1' & O"214",
    8#3176# => '1' & O"161",
    8#3177# => '1' & O"071",
    8#3200# => '1' & O"014",
    8#3201# => '1' & O"165",
    8#3202# => '0' & O"214",
    8#3203# => '1' & O"030",
    8#3204# => '0' & O"614",
    8#3205# => '1' & O"161",
    8#3206# => '0' & O"414",
    8#3207# => '1' & O"161",
    8#3210# => '1' & O"161",
    8#3211# => '1' & O"456",
    8#3212# => '1' & O"116",
    8#3213# => '1' & O"514",
    8#3214# => '0' & O"530",
    8#3215# => '1' & O"757",
    8#3216# => '0' & O"614",
    8#3217# => '1' & O"030",
    8#3220# => '0' & O"630",
    8#3221# => '0' & O"530",
    8#3222# => '0' & O"230",
    8#3223# => '0' & O"430",
    8#3224# => '1' & O"130",
    8#3225# => '0' & O"124",
    8#3226# => '1' & O"553",
    8#3227# => '0' & O"060",
    8#3230# => '1' & O"356",
    8#3231# => '1' & O"742",
    8#3232# => '1' & O"220",
    8#3233# => '1' & O"620",
    8#3234# => '0' & O"416",
    8#3235# => '1' & O"226",
    8#3236# => '1' & O"056",
    8#3237# => '1' & O"207",
    8#3240# => '0' & O"776",
    8#3241# => '1' & O"416",
    8#3242# => '1' & O"203",
    8#3243# => '1' & O"616",
    8#3244# => '1' & O"620",
    8#3245# => '1' & O"620",
    8#3246# => '0' & O"512",
    8#3247# => '1' & O"620",
    8#3250# => '0' & O"742",
    8#3251# => '1' & O"516",
    8#3252# => '1' & O"243",
    8#3253# => '1' & O"716",
    8#3254# => '0' & O"416",
    8#3255# => '0' & O"034",
    8#3256# => '1' & O"122",
    8#3257# => '0' & O"054",
    8#3260# => '1' & O"247",
    8#3261# => '0' & O"267",
    8#3262# => '0' & O"742",
    8#3263# => '1' & O"426",
    8#3264# => '1' & O"313",
    8#3265# => '1' & O"626",
    8#3266# => '0' & O"426",
    8#3267# => '0' & O"034",
    8#3270# => '0' & O"054",
    8#3271# => '1' & O"317",
    8#3272# => '0' & O"267",
    8#3273# => '0' & O"034",
    8#3274# => '1' & O"626",
    8#3275# => '1' & O"557",
    8#3276# => '0' & O"620",
    8#3277# => '0' & O"572",
    8#3300# => '0' & O"572",
    8#3301# => '1' & O"352",
    8#3302# => '1' & O"536",
    8#3303# => '1' & O"176",
    8#3304# => '1' & O"433",
    8#3305# => '1' & O"620",
    8#3306# => '1' & O"006",
    8#3307# => '1' & O"453",
    8#3310# => '0' & O"376",
    8#3311# => '1' & O"456",
    8#3312# => '1' & O"416",
    8#3313# => '1' & O"620",
    8#3314# => '0' & O"316",
    8#3315# => '1' & O"314",
    8#3316# => '0' & O"730",
    8#3317# => '1' & O"030",
    8#3320# => '0' & O"530",
    8#3321# => '0' & O"330",
    8#3322# => '1' & O"130",
    8#3323# => '1' & O"030",
    8#3324# => '0' & O"130",
    8#3325# => '0' & O"630",
    8#3326# => '0' & O"330",
    8#3327# => '0' & O"530",
    8#3330# => '1' & O"220",
    8#3331# => '0' & O"060",
    8#3332# => '0' & O"620",
    8#3333# => '1' & O"612",
    8#3334# => '1' & O"573",
    8#3335# => '0' & O"542",
    8#3336# => '0' & O"776",
    8#3337# => '0' & O"054",
    8#3340# => '1' & O"357",
    8#3341# => '1' & O"652",
    8#3342# => '1' & O"352",
    8#3343# => '0' & O"142",
    8#3344# => '1' & O"633",
    8#3345# => '1' & O"316",
    8#3346# => '1' & O"116",
    8#3347# => '1' & O"052",
    8#3350# => '0' & O"312",
    8#3351# => '1' & O"414",
    8#3352# => '1' & O"273",
    8#3353# => '1' & O"620",
    8#3354# => '1' & O"222",
    8#3355# => '1' & O"222",
    8#3356# => '0' & O"576",
    8#3357# => '1' & O"663",
    8#3360# => '0' & O"722",
    8#3361# => '1' & O"422",
    8#3362# => '1' & O"062",
    8#3363# => '0' & O"216",
    8#3364# => '1' & O"576",
    8#3365# => '1' & O"673",
    8#3366# => '1' & O"662",
    8#3367# => '0' & O"650",
    8#3370# => '0' & O"036",
    8#3371# => '0' & O"007",
    8#3372# => '0' & O"416",
    8#3373# => '1' & O"662",
    8#3374# => '0' & O"450",
    8#3375# => '1' & O"222",
    8#3376# => '0' & O"576",
    8#3377# => '1' & O"076",
    8#3400# => '0' & O"000",
    8#3401# => '1' & O"476",
    8#3402# => '1' & O"776",
    8#3403# => '1' & O"126",
    8#3404# => '0' & O"422",
    8#3405# => '0' & O"113",
    8#3406# => '0' & O"650",
    8#3407# => '1' & O"231",
    8#3410# => '0' & O"420",
    8#3411# => '1' & O"731",
    8#3412# => '0' & O"056",
    8#3413# => '1' & O"231",
    8#3414# => '0' & O"616",
    8#3415# => '0' & O"413",
    8#3416# => '0' & O"572",
    8#3417# => '1' & O"364",
    8#3420# => '0' & O"707",
    8#3421# => '0' & O"776",
    8#3422# => '0' & O"456",
    8#3423# => '1' & O"131",
    8#3424# => '1' & O"542",
    8#3425# => '0' & O"107",
    8#3426# => '1' & O"462",
    8#3427# => '1' & O"636",
    8#3430# => '0' & O"007",
    8#3431# => '0' & O"714",
    8#3432# => '0' & O"665",
    8#3433# => '1' & O"014",
    8#3434# => '1' & O"165",
    8#3435# => '1' & O"114",
    8#3436# => '1' & O"161",
    8#3437# => '1' & O"771",
    8#3440# => '1' & O"214",
    8#3441# => '1' & O"161",
    8#3442# => '0' & O"765",
    8#3443# => '1' & O"314",
    8#3444# => '1' & O"161",
    8#3445# => '1' & O"575",
    8#3446# => '1' & O"161",
    8#3447# => '1' & O"345",
    8#3450# => '1' & O"161",
    8#3451# => '1' & O"731",
    8#3452# => '1' & O"656",
    8#3453# => '0' & O"516",
    8#3454# => '0' & O"032",
    8#3455# => '0' & O"277",
    8#3456# => '0' & O"516",
    8#3457# => '1' & O"456",
    8#3460# => '0' & O"034",
    8#3461# => '0' & O"416",
    8#3462# => '0' & O"154",
    8#3463# => '0' & O"303",
    8#3464# => '1' & O"656",
    8#3465# => '0' & O"676",
    8#3466# => '0' & O"343",
    8#3467# => '0' & O"346",
    8#3470# => '0' & O"752",
    8#3471# => '1' & O"314",
    8#3472# => '1' & O"425",
    8#3473# => '1' & O"124",
    8#3474# => '0' & O"033",
    8#3475# => '0' & O"524",
    8#3476# => '1' & O"123",
    8#3477# => '1' & O"731",
    8#3500# => '1' & O"235",
    8#3501# => '1' & O"123",
    8#3502# => '1' & O"731",
    8#3503# => '1' & O"661",
    8#3504# => '1' & O"345",
    8#3505# => '1' & O"314",
    8#3506# => '1' & O"155",
    8#3507# => '1' & O"575",
    8#3510# => '1' & O"214",
    8#3511# => '1' & O"155",
    8#3512# => '0' & O"765",
    8#3513# => '1' & O"114",
    8#3514# => '1' & O"155",
    8#3515# => '1' & O"771",
    8#3516# => '1' & O"014",
    8#3517# => '1' & O"155",
    8#3520# => '1' & O"155",
    8#3521# => '1' & O"155",
    8#3522# => '0' & O"614",
    8#3523# => '1' & O"362",
    8#3524# => '1' & O"514",
    8#3525# => '1' & O"056",
    8#3526# => '1' & O"656",
    8#3527# => '0' & O"630",
    8#3530# => '1' & O"073",
    8#3531# => '0' & O"224",
    8#3532# => '0' & O"573",
    8#3533# => '1' & O"752",
    8#3534# => '1' & O"172",
    8#3535# => '1' & O"413",
    8#3536# => '1' & O"426",
    8#3537# => '0' & O"547",
    8#3540# => '1' & O"626",
    8#3541# => '0' & O"416",
    8#3542# => '0' & O"552",
    8#3543# => '0' & O"563",
    8#3544# => '1' & O"316",
    8#3545# => '0' & O"322",
    8#3546# => '1' & O"652",
    8#3547# => '0' & O"676",
    8#3550# => '0' & O"663",
    8#3551# => '1' & O"456",
    8#3552# => '1' & O"416",
    8#3553# => '0' & O"356",
    8#3554# => '1' & O"316",
    8#3555# => '1' & O"056",
    8#3556# => '0' & O"316",
    8#3557# => '0' & O"546",
    8#3560# => '0' & O"224",
    8#3561# => '0' & O"733",
    8#3562# => '0' & O"430",
    8#3563# => '0' & O"746",
    8#3564# => '0' & O"747",
    8#3565# => '0' & O"630",
    8#3566# => '0' & O"154",
    8#3567# => '0' & O"727",
    8#3570# => '1' & O"116",
    8#3571# => '1' & O"116",
    8#3572# => '0' & O"224",
    8#3573# => '1' & O"123",
    8#3574# => '0' & O"060",
    8#3575# => '0' & O"714",
    8#3576# => '0' & O"330",
    8#3577# => '0' & O"330",
    8#3600# => '0' & O"030",
    8#3601# => '1' & O"030",
    8#3602# => '0' & O"530",
    8#3603# => '0' & O"030",
    8#3604# => '1' & O"130",
    8#3605# => '1' & O"653",
    8#3606# => '1' & O"131",
    8#3607# => '1' & O"742",
    8#3610# => '0' & O"456",
    8#3611# => '0' & O"576",
    8#3612# => '1' & O"033",
    8#3613# => '1' & O"322",
    8#3614# => '1' & O"656",
    8#3615# => '0' & O"426",
    8#3616# => '1' & O"656",
    8#3617# => '1' & O"576",
    8#3620# => '1' & O"043",
    8#3621# => '1' & O"456",
    8#3622# => '1' & O"742",
    8#3623# => '1' & O"461",
    8#3624# => '1' & O"420",
    8#3625# => '1' & O"322",
    8#3626# => '1' & O"576",
    8#3627# => '1' & O"127",
    8#3630# => '1' & O"376",
    8#3631# => '1' & O"616",
    8#3632# => '0' & O"060",
    8#3633# => '1' & O"420",
    8#3634# => '1' & O"316",
    8#3635# => '1' & O"056",
    8#3636# => '1' & O"203",
    8#3637# => '1' & O"616",
    8#3640# => '0' & O"576",
    8#3641# => '1' & O"177",
    8#3642# => '1' & O"656",
    8#3643# => '0' & O"426",
    8#3644# => '1' & O"656",
    8#3645# => '0' & O"667",
    8#3646# => '0' & O"314",
    8#3647# => '0' & O"712",
    8#3650# => '0' & O"536",
    8#3651# => '1' & O"257",
    8#3652# => '0' & O"276",
    8#3653# => '1' & O"446",
    8#3654# => '1' & O"356",
    8#3655# => '1' & O"454",
    8#3656# => '1' & O"427",
    8#3657# => '0' & O"146",
    8#3660# => '1' & O"333",
    8#3661# => '0' & O"322",
    8#3662# => '0' & O"562",
    8#3663# => '0' & O"332",
    8#3664# => '1' & O"557",
    8#3665# => '0' & O"000",
    8#3666# => '1' & O"062",
    8#3667# => '1' & O"646",
    8#3670# => '1' & O"420",
    8#3671# => '1' & O"244",
    8#3672# => '0' & O"630",
    8#3673# => '1' & O"130",
    8#3674# => '0' & O"330",
    8#3675# => '0' & O"130",
    8#3676# => '0' & O"430",
    8#3677# => '0' & O"730",
    8#3700# => '0' & O"130",
    8#3701# => '1' & O"633",
    8#3702# => '1' & O"746",
    8#3703# => '0' & O"623",
    8#3704# => '1' & O"616",
    8#3705# => '0' & O"542",
    8#3706# => '1' & O"423",
    8#3707# => '1' & O"316",
    8#3710# => '0' & O"074",
    8#3711# => '1' & O"554",
    8#3712# => '1' & O"427",
    8#3713# => '0' & O"752",
    8#3714# => '1' & O"376",
    8#3715# => '1' & O"414",
    8#3716# => '0' & O"056",
    8#3717# => '1' & O"142",
    8#3720# => '1' & O"533",
    8#3721# => '0' & O"416",
    8#3722# => '0' & O"552",
    8#3723# => '1' & O"156",
    8#3724# => '1' & O"477",
    8#3725# => '0' & O"316",
    8#3726# => '0' & O"452",
    8#3727# => '1' & O"616",
    8#3730# => '1' & O"176",
    8#3731# => '1' & O"437",
    8#3732# => '1' & O"646",
    8#3733# => '0' & O"616",
    8#3734# => '0' & O"056",
    8#3735# => '1' & O"414",
    8#3736# => '0' & O"753",
    8#3737# => '1' & O"114",
    8#3740# => '0' & O"330",
    8#3741# => '0' & O"130",
    8#3742# => '0' & O"030",
    8#3743# => '0' & O"130",
    8#3744# => '0' & O"730",
    8#3745# => '1' & O"130",
    8#3746# => '1' & O"030",
    8#3747# => '0' & O"030",
    8#3750# => '0' & O"530",
    8#3751# => '0' & O"530",
    8#3752# => '0' & O"330",
    8#3753# => '1' & O"567",
    8#3754# => '1' & O"656",
    8#3755# => '0' & O"456",
    8#3756# => '0' & O"606",
    8#3757# => '1' & O"272",
    8#3760# => '0' & O"573",
    8#3761# => '0' & O"772",
    8#3762# => '1' & O"316",
    8#3763# => '0' & O"752",
    8#3764# => '1' & O"713",
    8#3765# => '0' & O"637",
    8#3766# => '0' & O"316",
    8#3767# => '1' & O"414",
    8#3770# => '0' & O"230",
    8#3771# => '0' & O"330",
    8#3772# => '0' & O"030",
    8#3773# => '0' & O"230",
    8#3774# => '0' & O"530",
    8#3775# => '1' & O"007",
    8#3776# => '0' & O"514",
    8#3777# => '0' & O"773",
    8#4000# => '0' & O"220",
    8#4001# => '0' & O"742",
    8#4002# => '0' & O"742",
    8#4003# => '0' & O"742",
    8#4004# => '0' & O"742",
    8#4005# => '0' & O"000",
    8#4006# => '0' & O"742",
    8#4007# => '0' & O"413",
    8#4010# => '0' & O"250",
    8#4011# => '0' & O"143",
    8#4012# => '0' & O"742",
    8#4013# => '0' & O"742",
    8#4014# => '0' & O"742",
    8#4015# => '0' & O"000",
    8#4016# => '0' & O"742",
    8#4017# => '0' & O"403",
    8#4020# => '0' & O"364",
    8#4021# => '1' & O"617",
    8#4022# => '0' & O"742",
    8#4023# => '0' & O"742",
    8#4024# => '0' & O"742",
    8#4025# => '0' & O"153",
    8#4026# => '1' & O"030",
    8#4027# => '0' & O"403",
    8#4030# => '0' & O"364",
    8#4031# => '0' & O"617",
    8#4032# => '0' & O"742",
    8#4033# => '0' & O"742",
    8#4034# => '0' & O"742",
    8#4035# => '0' & O"417",
    8#4036# => '1' & O"030",
    8#4037# => '0' & O"407",
    8#4040# => '0' & O"000",
    8#4041# => '0' & O"742",
    8#4042# => '0' & O"007",
    8#4043# => '0' & O"207",
    8#4044# => '0' & O"417",
    8#4045# => '0' & O"000",
    8#4046# => '1' & O"030",
    8#4047# => '0' & O"413",
    8#4050# => '0' & O"504",
    8#4051# => '0' & O"003",
    8#4052# => '0' & O"742",
    8#4053# => '0' & O"742",
    8#4054# => '0' & O"742",
    8#4055# => '0' & O"000",
    8#4056# => '0' & O"742",
    8#4057# => '0' & O"407",
    8#4060# => '1' & O"306",
    8#4061# => '1' & O"061",
    8#4062# => '0' & O"742",
    8#4063# => '0' & O"742",
    8#4064# => '0' & O"742",
    8#4065# => '0' & O"113",
    8#4066# => '1' & O"030",
    8#4067# => '0' & O"377",
    8#4070# => '0' & O"742",
    8#4071# => '0' & O"000",
    8#4072# => '0' & O"742",
    8#4073# => '0' & O"742",
    8#4074# => '0' & O"000",
    8#4075# => '0' & O"000",
    8#4076# => '0' & O"742",
    8#4077# => '0' & O"772",
    8#4100# => '0' & O"772",
    8#4101# => '0' & O"772",
    8#4102# => '0' & O"772",
    8#4103# => '0' & O"114",
    8#4104# => '0' & O"324",
    8#4105# => '1' & O"273",
    8#4106# => '0' & O"612",
    8#4107# => '0' & O"250",
    8#4110# => '0' & O"676",
    8#4111# => '1' & O"643",
    8#4112# => '0' & O"576",
    8#4113# => '0' & O"676",
    8#4114# => '0' & O"103",
    8#4115# => '0' & O"250",
    8#4116# => '0' & O"312",
    8#4117# => '0' & O"530",
    8#4120# => '0' & O"112",
    8#4121# => '1' & O"637",
    8#4122# => '1' & O"712",
    8#4123# => '0' & O"512",
    8#4124# => '1' & O"326",
    8#4125# => '0' & O"412",
    8#4126# => '0' & O"416",
    8#4127# => '0' & O"612",
    8#4130# => '0' & O"316",
    8#4131# => '0' & O"566",
    8#4132# => '0' & O"542",
    8#4133# => '0' & O"000",
    8#4134# => '1' & O"572",
    8#4135# => '0' & O"514",
    8#4136# => '0' & O"030",
    8#4137# => '0' & O"230",
    8#4140# => '1' & O"376",
    8#4141# => '1' & O"056",
    8#4142# => '1' & O"314",
    8#4143# => '0' & O"250",
    8#4144# => '0' & O"302",
    8#4145# => '0' & O"044",
    8#4146# => '0' & O"034",
    8#4147# => '1' & O"354",
    8#4150# => '0' & O"633",
    8#4151# => '1' & O"050",
    8#4152# => '0' & O"642",
    8#4153# => '0' & O"737",
    8#4154# => '0' & O"524",
    8#4155# => '0' & O"677",
    8#4156# => '1' & O"103",
    8#4157# => '0' & O"250",
    8#4160# => '1' & O"124",
    8#4161# => '0' & O"727",
    8#4162# => '0' & O"114",
    8#4163# => '0' & O"312",
    8#4164# => '0' & O"320",
    8#4165# => '1' & O"056",
    8#4166# => '0' & O"713",
    8#4167# => '0' & O"050",
    8#4170# => '0' & O"024",
    8#4171# => '0' & O"757",
    8#4172# => '0' & O"627",
    8#4173# => '0' & O"302",
    8#4174# => '0' & O"742",
    8#4175# => '0' & O"344",
    8#4176# => '1' & O"344",
    8#4177# => '1' & O"000",
    8#4200# => '0' & O"524",
    8#4201# => '1' & O"647",
    8#4202# => '0' & O"034",
    8#4203# => '1' & O"354",
    8#4204# => '1' & O"003",
    8#4205# => '0' & O"776",
    8#4206# => '1' & O"003",
    8#4207# => '0' & O"737",
    8#4210# => '1' & O"722",
    8#4211# => '1' & O"522",
    8#4212# => '1' & O"607",
    8#4213# => '1' & O"514",
    8#4214# => '1' & O"752",
    8#4215# => '0' & O"303",
    8#4216# => '1' & O"333",
    8#4217# => '0' & O"000",
    8#4220# => '0' & O"336",
    8#4221# => '0' & O"250",
    8#4222# => '0' & O"064",
    8#4223# => '0' & O"704",
    8#4224# => '1' & O"124",
    8#4225# => '1' & O"143",
    8#4226# => '1' & O"044",
    8#4227# => '0' & O"613",
    8#4230# => '0' & O"616",
    8#4231# => '1' & O"250",
    8#4232# => '0' & O"456",
    8#4233# => '1' & O"104",
    8#4234# => '1' & O"014",
    8#4235# => '0' & O"034",
    8#4236# => '1' & O"116",
    8#4237# => '0' & O"154",
    8#4240# => '1' & O"167",
    8#4241# => '0' & O"142",
    8#4242# => '1' & O"317",
    8#4243# => '1' & O"172",
    8#4244# => '1' & O"043",
    8#4245# => '1' & O"142",
    8#4246# => '1' & O"607",
    8#4247# => '1' & O"514",
    8#4250# => '0' & O"034",
    8#4251# => '1' & O"552",
    8#4252# => '1' & O"243",
    8#4253# => '1' & O"333",
    8#4254# => '1' & O"144",
    8#4255# => '1' & O"133",
    8#4256# => '1' & O"112",
    8#4257# => '0' & O"220",
    8#4260# => '1' & O"024",
    8#4261# => '0' & O"743",
    8#4262# => '1' & O"103",
    8#4263# => '1' & O"144",
    8#4264# => '0' & O"302",
    8#4265# => '1' & O"414",
    8#4266# => '0' & O"326",
    8#4267# => '0' & O"742",
    8#4270# => '0' & O"742",
    8#4271# => '0' & O"034",
    8#4272# => '0' & O"254",
    8#4273# => '1' & O"427",
    8#4274# => '0' & O"312",
    8#4275# => '1' & O"656",
    8#4276# => '1' & O"124",
    8#4277# => '1' & O"543",
    8#4300# => '1' & O"552",
    8#4301# => '1' & O"541",
    8#4302# => '0' & O"742",
    8#4303# => '1' & O"763",
    8#4304# => '1' & O"463",
    8#4305# => '0' & O"552",
    8#4306# => '1' & O"347",
    8#4307# => '0' & O"322",
    8#4310# => '0' & O"562",
    8#4311# => '1' & O"656",
    8#4312# => '1' & O"242",
    8#4313# => '1' & O"763",
    8#4314# => '0' & O"074",
    8#4315# => '1' & O"554",
    8#4316# => '1' & O"413",
    8#4317# => '0' & O"034",
    8#4320# => '0' & O"306",
    8#4321# => '0' & O"742",
    8#4322# => '1' & O"124",
    8#4323# => '1' & O"533",
    8#4324# => '1' & O"326",
    8#4325# => '1' & O"552",
    8#4326# => '0' & O"752",
    8#4327# => '1' & O"752",
    8#4330# => '0' & O"772",
    8#4331# => '1' & O"573",
    8#4332# => '0' & O"252",
    8#4333# => '1' & O"656",
    8#4334# => '1' & O"056",
    8#4335# => '1' & O"263",
    8#4336# => '0' & O"572",
    8#4337# => '0' & O"672",
    8#4340# => '1' & O"557",
    8#4341# => '1' & O"456",
    8#4342# => '1' & O"250",
    8#4343# => '1' & O"014",
    8#4344# => '0' & O"130",
    8#4345# => '1' & O"130",
    8#4346# => '1' & O"153",
    8#4347# => '0' & O"250",
    8#4350# => '0' & O"220",
    8#4351# => '1' & O"324",
    8#4352# => '1' & O"667",
    8#4353# => '1' & O"711",
    8#4354# => '0' & O"620",
    8#4355# => '0' & O"324",
    8#4356# => '1' & O"303",
    8#4357# => '1' & O"024",
    8#4360# => '1' & O"747",
    8#4361# => '0' & O"743",
    8#4362# => '0' & O"336",
    8#4363# => '0' & O"250",
    8#4364# => '1' & O"124",
    8#4365# => '1' & O"737",
    8#4366# => '0' & O"060",
    8#4367# => '1' & O"056",
    8#4370# => '0' & O"060",
    8#4371# => '1' & O"711",
    8#4372# => '1' & O"064",
    8#4373# => '1' & O"220",
    8#4374# => '1' & O"124",
    8#4375# => '1' & O"537",
    8#4376# => '0' & O"332",
    8#4377# => '1' & O"541",
    8#4400# => '0' & O"000",
    8#4401# => '0' & O"250",
    8#4402# => '0' & O"324",
    8#4403# => '0' & O"177",
    8#4404# => '0' & O"616",
    8#4405# => '0' & O"316",
    8#4406# => '0' & O"746",
    8#4407# => '0' & O"414",
    8#4410# => '0' & O"524",
    8#4411# => '0' & O"077",
    8#4412# => '0' & O"544",
    8#4413# => '1' & O"722",
    8#4414# => '1' & O"656",
    8#4415# => '0' & O"250",
    8#4416# => '0' & O"367",
    8#4417# => '1' & O"522",
    8#4420# => '0' & O"061",
    8#4421# => '0' & O"114",
    8#4422# => '1' & O"656",
    8#4423# => '0' & O"642",
    8#4424# => '0' & O"137",
    8#4425# => '0' & O"352",
    8#4426# => '0' & O"332",
    8#4427# => '0' & O"612",
    8#4430# => '0' & O"477",
    8#4431# => '1' & O"116",
    8#4432# => '0' & O"034",
    8#4433# => '1' & O"267",
    8#4434# => '1' & O"116",
    8#4435# => '0' & O"034",
    8#4436# => '0' & O"377",
    8#4437# => '0' & O"524",
    8#4440# => '1' & O"207",
    8#4441# => '0' & O"544",
    8#4442# => '1' & O"167",
    8#4443# => '1' & O"522",
    8#4444# => '1' & O"567",
    8#4445# => '1' & O"414",
    8#4446# => '0' & O"322",
    8#4447# => '0' & O"562",
    8#4450# => '0' & O"414",
    8#4451# => '1' & O"317",
    8#4452# => '0' & O"000",
    8#4453# => '0' & O"312",
    8#4454# => '0' & O"154",
    8#4455# => '0' & O"317",
    8#4456# => '0' & O"652",
    8#4457# => '0' & O"337",
    8#4460# => '0' & O"552",
    8#4461# => '0' & O"074",
    8#4462# => '0' & O"273",
    8#4463# => '0' & O"752",
    8#4464# => '0' & O"416",
    8#4465# => '0' & O"034",
    8#4466# => '0' & O"263",
    8#4467# => '1' & O"370",
    8#4470# => '1' & O"642",
    8#4471# => '0' & O"034",
    8#4472# => '1' & O"642",
    8#4473# => '1' & O"360",
    8#4474# => '1' & O"775",
    8#4475# => '1' & O"711",
    8#4476# => '1' & O"370",
    8#4477# => '0' & O"154",
    8#4500# => '0' & O"163",
    8#4501# => '0' & O"747",
    8#4502# => '0' & O"612",
    8#4503# => '0' & O"312",
    8#4504# => '0' & O"114",
    8#4505# => '0' & O"530",
    8#4506# => '1' & O"372",
    8#4507# => '1' & O"512",
    8#4510# => '0' & O"473",
    8#4511# => '1' & O"712",
    8#4512# => '1' & O"112",
    8#4513# => '0' & O"102",
    8#4514# => '0' & O"107",
    8#4515# => '0' & O"477",
    8#4516# => '1' & O"572",
    8#4517# => '1' & O"250",
    8#4520# => '0' & O"606",
    8#4521# => '0' & O"406",
    8#4522# => '0' & O"316",
    8#4523# => '0' & O"566",
    8#4524# => '0' & O"752",
    8#4525# => '1' & O"324",
    8#4526# => '0' & O"543",
    8#4527# => '0' & O"312",
    8#4530# => '0' & O"552",
    8#4531# => '0' & O"250",
    8#4532# => '0' & O"336",
    8#4533# => '0' & O"250",
    8#4534# => '0' & O"020",
    8#4535# => '0' & O"336",
    8#4536# => '0' & O"644",
    8#4537# => '0' & O"444",
    8#4540# => '0' & O"244",
    8#4541# => '0' & O"144",
    8#4542# => '0' & O"060",
    8#4543# => '0' & O"336",
    8#4544# => '0' & O"776",
    8#4545# => '0' & O"776",
    8#4546# => '0' & O"250",
    8#4547# => '0' & O"324",
    8#4550# => '0' & O"763",
    8#4551# => '1' & O"250",
    8#4552# => '0' & O"746",
    8#4553# => '0' & O"606",
    8#4554# => '0' & O"414",
    8#4555# => '1' & O"242",
    8#4556# => '0' & O"713",
    8#4557# => '0' & O"030",
    8#4560# => '0' & O"030",
    8#4561# => '1' & O"653",
    8#4562# => '0' & O"406",
    8#4563# => '0' & O"316",
    8#4564# => '0' & O"556",
    8#4565# => '0' & O"332",
    8#4566# => '1' & O"372",
    8#4567# => '1' & O"572",
    8#4570# => '0' & O"561",
    8#4571# => '1' & O"324",
    8#4572# => '1' & O"703",
    8#4573# => '0' & O"413",
    8#4574# => '0' & O"601",
    8#4575# => '1' & O"124",
    8#4576# => '1' & O"003",
    8#4577# => '1' & O"007",
    8#4600# => '1' & O"056",
    8#4601# => '0' & O"250",
    8#4602# => '1' & O"414",
    8#4603# => '1' & O"024",
    8#4604# => '1' & O"067",
    8#4605# => '1' & O"314",
    8#4606# => '0' & O"044",
    8#4607# => '0' & O"024",
    8#4610# => '1' & O"137",
    8#4611# => '0' & O"142",
    8#4612# => '1' & O"143",
    8#4613# => '1' & O"414",
    8#4614# => '1' & O"117",
    8#4615# => '0' & O"642",
    8#4616# => '1' & O"117",
    8#4617# => '0' & O"746",
    8#4620# => '0' & O"742",
    8#4621# => '0' & O"542",
    8#4622# => '1' & O"027",
    8#4623# => '0' & O"302",
    8#4624# => '0' & O"250",
    8#4625# => '0' & O"164",
    8#4626# => '1' & O"123",
    8#4627# => '0' & O"302",
    8#4630# => '0' & O"050",
    8#4631# => '0' & O"250",
    8#4632# => '1' & O"124",
    8#4633# => '1' & O"233",
    8#4634# => '1' & O"237",
    8#4635# => '1' & O"414",
    8#4636# => '1' & O"130",
    8#4637# => '0' & O"250",
    8#4640# => '1' & O"237",
    8#4641# => '0' & O"565",
    8#4642# => '0' & O"414",
    8#4643# => '0' & O"322",
    8#4644# => '0' & O"250",
    8#4645# => '0' & O"767",
    8#4646# => '1' & O"056",
    8#4647# => '1' & O"711",
    8#4650# => '1' & O"324",
    8#4651# => '1' & O"263",
    8#4652# => '1' & O"064",
    8#4653# => '0' & O"037",
    8#4654# => '1' & O"370",
    8#4655# => '0' & O"154",
    8#4656# => '0' & O"147",
    8#4657# => '1' & O"775",
    8#4660# => '0' & O"114",
    8#4661# => '1' & O"064",
    8#4662# => '0' & O"103",
    8#4663# => '1' & O"662",
    8#4664# => '0' & O"622",
    8#4665# => '1' & O"714",
    8#4666# => '0' & O"034",
    8#4667# => '0' & O"034",
    8#4670# => '0' & O"746",
    8#4671# => '1' & O"333",
    8#4672# => '1' & O"116",
    8#4673# => '0' & O"776",
    8#4674# => '0' & O"776",
    8#4675# => '1' & O"116",
    8#4676# => '0' & O"312",
    8#4677# => '0' & O"752",
    8#4700# => '1' & O"160",
    8#4701# => '0' & O"312",
    8#4702# => '0' & O"552",
    8#4703# => '0' & O"552",
    8#4704# => '0' & O"552",
    8#4705# => '1' & O"656",
    8#4706# => '0' & O"412",
    8#4707# => '1' & O"372",
    8#4710# => '0' & O"416",
    8#4711# => '0' & O"416",
    8#4712# => '1' & O"656",
    8#4713# => '0' & O"576",
    8#4714# => '0' & O"576",
    8#4715# => '0' & O"576",
    8#4716# => '1' & O"523",
    8#4717# => '1' & O"746",
    8#4720# => '0' & O"250",
    8#4721# => '1' & O"656",
    8#4722# => '0' & O"250",
    8#4723# => '0' & O"060",
    8#4724# => '1' & O"706",
    8#4725# => '1' & O"467",
    8#4726# => '1' & O"662",
    8#4727# => '0' & O"314",
    8#4730# => '0' & O"730",
    8#4731# => '0' & O"414",
    8#4732# => '1' & O"546",
    8#4733# => '0' & O"776",
    8#4734# => '0' & O"776",
    8#4735# => '0' & O"776",
    8#4736# => '0' & O"217",
    8#4737# => '1' & O"656",
    8#4740# => '0' & O"322",
    8#4741# => '0' & O"606",
    8#4742# => '1' & O"733",
    8#4743# => '0' & O"250",
    8#4744# => '1' & O"172",
    8#4745# => '1' & O"643",
    8#4746# => '0' & O"412",
    8#4747# => '1' & O"316",
    8#4750# => '0' & O"250",
    8#4751# => '0' & O"746",
    8#4752# => '0' & O"250",
    8#4753# => '1' & O"312",
    8#4754# => '1' & O"711",
    8#4755# => '1' & O"324",
    8#4756# => '0' & O"257",
    8#4757# => '0' & O"367",
    8#4760# => '1' & O"775",
    8#4761# => '0' & O"413",
    8#4762# => '1' & O"344",
    8#4763# => '0' & O"250",
    8#4764# => '1' & O"656",
    8#4765# => '0' & O"250",
    8#4766# => '0' & O"316",
    8#4767# => '0' & O"414",
    8#4770# => '1' & O"662",
    8#4771# => '0' & O"146",
    8#4772# => '1' & O"533",
    8#4773# => '1' & O"662",
    8#4774# => '1' & O"304",
    8#4775# => '1' & O"503",
    8#4776# => '0' & O"000",
    8#4777# => '0' & O"420",
    8#5000# => '0' & O"250",
    8#5001# => '0' & O"514",
    8#5002# => '0' & O"542",
    8#5003# => '0' & O"364",
    8#5004# => '1' & O"513",
    8#5005# => '0' & O"752",
    8#5006# => '1' & O"316",
    8#5007# => '0' & O"056",
    8#5010# => '0' & O"452",
    8#5011# => '1' & O"616",
    8#5012# => '1' & O"176",
    8#5013# => '0' & O"027",
    8#5014# => '1' & O"623",
    8#5015# => '0' & O"032",
    8#5016# => '1' & O"463",
    8#5017# => '1' & O"517",
    8#5020# => '1' & O"552",
    8#5021# => '0' & O"637",
    8#5022# => '0' & O"430",
    8#5023# => '0' & O"530",
    8#5024# => '0' & O"330",
    8#5025# => '0' & O"530",
    8#5026# => '1' & O"130",
    8#5027# => '0' & O"230",
    8#5030# => '0' & O"330",
    8#5031# => '0' & O"730",
    8#5032# => '0' & O"343",
    8#5033# => '1' & O"552",
    8#5034# => '0' & O"103",
    8#5035# => '0' & O"130",
    8#5036# => '0' & O"030",
    8#5037# => '0' & O"530",
    8#5040# => '0' & O"530",
    8#5041# => '0' & O"030",
    8#5042# => '0' & O"530",
    8#5043# => '0' & O"530",
    8#5044# => '1' & O"030",
    8#5045# => '0' & O"530",
    8#5046# => '0' & O"330",
    8#5047# => '0' & O"014",
    8#5050# => '0' & O"330",
    8#5051# => '0' & O"347",
    8#5052# => '1' & O"414",
    8#5053# => '1' & O"552",
    8#5054# => '0' & O"157",
    8#5055# => '0' & O"130",
    8#5056# => '0' & O"730",
    8#5057# => '0' & O"430",
    8#5060# => '0' & O"530",
    8#5061# => '0' & O"330",
    8#5062# => '0' & O"230",
    8#5063# => '1' & O"130",
    8#5064# => '0' & O"230",
    8#5065# => '0' & O"530",
    8#5066# => '0' & O"230",
    8#5067# => '0' & O"552",
    8#5070# => '0' & O"552",
    8#5071# => '1' & O"064",
    8#5072# => '1' & O"707",
    8#5073# => '1' & O"552",
    8#5074# => '0' & O"413",
    8#5075# => '0' & O"230",
    8#5076# => '0' & O"530",
    8#5077# => '0' & O"430",
    8#5100# => '0' & O"752",
    8#5101# => '0' & O"347",
    8#5102# => '1' & O"552",
    8#5103# => '1' & O"727",
    8#5104# => '0' & O"330",
    8#5105# => '0' & O"030",
    8#5106# => '0' & O"430",
    8#5107# => '1' & O"030",
    8#5110# => '0' & O"343",
    8#5111# => '1' & O"552",
    8#5112# => '0' & O"357",
    8#5113# => '0' & O"504",
    8#5114# => '0' & O"347",
    8#5115# => '0' & O"542",
    8#5116# => '0' & O"642",
    8#5117# => '0' & O"523",
    8#5120# => '1' & O"130",
    8#5121# => '0' & O"523",
    8#5122# => '1' & O"004",
    8#5123# => '0' & O"130",
    8#5124# => '0' & O"364",
    8#5125# => '1' & O"013",
    8#5126# => '0' & O"000",
    8#5127# => '0' & O"000",
    8#5130# => '1' & O"414",
    8#5131# => '0' & O"176",
    8#5132# => '0' & O"777",
    8#5133# => '0' & O"172",
    8#5134# => '0' & O"777",
    8#5135# => '0' & O"616",
    8#5136# => '0' & O"456",
    8#5137# => '0' & O"426",
    8#5140# => '1' & O"162",
    8#5141# => '1' & O"043",
    8#5142# => '1' & O"752",
    8#5143# => '0' & O"112",
    8#5144# => '1' & O"057",
    8#5145# => '0' & O"772",
    8#5146# => '1' & O"263",
    8#5147# => '1' & O"552",
    8#5150# => '0' & O"447",
    8#5151# => '0' & O"430",
    8#5152# => '0' & O"430",
    8#5153# => '0' & O"430",
    8#5154# => '1' & O"030",
    8#5155# => '0' & O"230",
    8#5156# => '0' & O"230",
    8#5157# => '0' & O"130",
    8#5160# => '0' & O"630",
    8#5161# => '0' & O"130",
    8#5162# => '0' & O"530",
    8#5163# => '0' & O"347",
    8#5164# => '0' & O"630",
    8#5165# => '0' & O"164",
    8#5166# => '1' & O"107",
    8#5167# => '0' & O"000",
    8#5170# => '0' & O"000",
    8#5171# => '0' & O"000",
    8#5172# => '0' & O"000",
    8#5173# => '0' & O"250",
    8#5174# => '1' & O"014",
    8#5175# => '0' & O"030",
    8#5176# => '0' & O"723",
    8#5177# => '1' & O"064",
    8#5200# => '0' & O"503",
    8#5201# => '0' & O"016",
    8#5202# => '1' & O"477",
    8#5203# => '1' & O"414",
    8#5204# => '0' & O"212",
    8#5205# => '1' & O"443",
    8#5206# => '1' & O"064",
    8#5207# => '0' & O"020",
    8#5210# => '1' & O"552",
    8#5211# => '0' & O"573",
    8#5212# => '0' & O"777",
    8#5213# => '0' & O"316",
    8#5214# => '0' & O"742",
    8#5215# => '1' & O"116",
    8#5216# => '0' & O"776",
    8#5217# => '1' & O"056",
    8#5220# => '0' & O"002",
    8#5221# => '1' & O"123",
    8#5222# => '1' & O"222",
    8#5223# => '0' & O"752",
    8#5224# => '1' & O"356",
    8#5225# => '1' & O"502",
    8#5226# => '1' & O"153",
    8#5227# => '0' & O"416",
    8#5230# => '1' & O"616",
    8#5231# => '1' & O"143",
    8#5232# => '1' & O"536",
    8#5233# => '1' & O"207",
    8#5234# => '1' & O"322",
    8#5235# => '1' & O"756",
    8#5236# => '0' & O"752",
    8#5237# => '1' & O"616",
    8#5240# => '1' & O"177",
    8#5241# => '1' & O"462",
    8#5242# => '0' & O"542",
    8#5243# => '1' & O"103",
    8#5244# => '0' & O"576",
    8#5245# => '1' & O"103",
    8#5246# => '0' & O"416",
    8#5247# => '0' & O"452",
    8#5250# => '1' & O"622",
    8#5251# => '0' & O"326",
    8#5252# => '1' & O"716",
    8#5253# => '1' & O"666",
    8#5254# => '1' & O"064",
    8#5255# => '1' & O"037",
    8#5256# => '1' & O"122",
    8#5257# => '0' & O"722",
    8#5260# => '0' & O"622",
    8#5261# => '1' & O"122",
    8#5262# => '1' & O"262",
    8#5263# => '1' & O"262",
    8#5264# => '0' & O"522",
    8#5265# => '0' & O"424",
    8#5266# => '1' & O"417",
    8#5267# => '0' & O"060",
    8#5270# => '1' & O"552",
    8#5271# => '0' & O"253",
    8#5272# => '0' & O"704",
    8#5273# => '1' & O"007",
    8#5274# => '1' & O"414",
    8#5275# => '0' & O"642",
    8#5276# => '0' & O"513",
    8#5277# => '1' & O"024",
    8#5300# => '0' & O"467",
    8#5301# => '1' & O"044",
    8#5302# => '0' & O"523",
    8#5303# => '1' & O"722",
    8#5304# => '1' & O"122",
    8#5305# => '0' & O"162",
    8#5306# => '1' & O"417",
    8#5307# => '0' & O"060",
    8#5310# => '0' & O"752",
    8#5311# => '0' & O"752",
    8#5312# => '0' & O"172",
    8#5313# => '0' & O"067",
    8#5314# => '0' & O"034",
    8#5315# => '0' & O"054",
    8#5316# => '1' & O"507",
    8#5317# => '0' & O"216",
    8#5320# => '1' & O"033",
    8#5321# => '0' & O"552",
    8#5322# => '1' & O"463",
    8#5323# => '0' & O"316",
    8#5324# => '0' & O"206",
    8#5325# => '0' & O"424",
    8#5326# => '1' & O"633",
    8#5327# => '0' & O"074",
    8#5330# => '0' & O"074",
    8#5331# => '1' & O"301",
    8#5332# => '0' & O"034",
    8#5333# => '0' & O"034",
    8#5334# => '1' & O"301",
    8#5335# => '0' & O"616",
    8#5336# => '0' & O"216",
    8#5337# => '1' & O"414",
    8#5340# => '1' & O"142",
    8#5341# => '1' & O"623",
    8#5342# => '0' & O"552",
    8#5343# => '0' & O"416",
    8#5344# => '1' & O"646",
    8#5345# => '1' & O"033",
    8#5346# => '1' & O"356",
    8#5347# => '1' & O"271",
    8#5350# => '0' & O"074",
    8#5351# => '0' & O"074",
    8#5352# => '1' & O"271",
    8#5353# => '0' & O"416",
    8#5354# => '0' & O"716",
    8#5355# => '1' & O"356",
    8#5356# => '0' & O"612",
    8#5357# => '1' & O"716",
    8#5360# => '0' & O"216",
    8#5361# => '1' & O"176",
    8#5362# => '0' & O"027",
    8#5363# => '1' & O"623",
    8#5364# => '0' & O"000",
    8#5365# => '0' & O"330",
    8#5366# => '0' & O"730",
    8#5367# => '1' & O"030",
    8#5370# => '0' & O"530",
    8#5371# => '0' & O"430",
    8#5372# => '0' & O"130",
    8#5373# => '0' & O"130",
    8#5374# => '0' & O"730",
    8#5375# => '1' & O"030",
    8#5376# => '0' & O"430",
    8#5377# => '0' & O"347",
    8#5400# => '0' & O"347",
    8#5401# => '1' & O"103",
    8#5402# => '0' & O"347",
    8#5403# => '0' & O"347",
    8#5404# => '0' & O"347",
    8#5405# => '0' & O"037",
    8#5406# => '0' & O"347",
    8#5407# => '0' & O"047",
    8#5410# => '0' & O"347",
    8#5411# => '0' & O"067",
    8#5412# => '0' & O"347",
    8#5413# => '0' & O"347",
    8#5414# => '0' & O"347",
    8#5415# => '0' & O"127",
    8#5416# => '0' & O"347",
    8#5417# => '0' & O"624",
    8#5420# => '0' & O"007",
    8#5421# => '0' & O"603",
    8#5422# => '0' & O"363",
    8#5423# => '0' & O"767",
    8#5424# => '0' & O"777",
    8#5425# => '0' & O"147",
    8#5426# => '0' & O"347",
    8#5427# => '1' & O"130",
    8#5430# => '1' & O"447",
    8#5431# => '0' & O"167",
    8#5432# => '1' & O"007",
    8#5433# => '1' & O"713",
    8#5434# => '1' & O"723",
    8#5435# => '0' & O"207",
    8#5436# => '0' & O"347",
    8#5437# => '1' & O"030",
    8#5440# => '1' & O"447",
    8#5441# => '0' & O"227",
    8#5442# => '1' & O"043",
    8#5443# => '0' & O"347",
    8#5444# => '1' & O"733",
    8#5445# => '0' & O"237",
    8#5446# => '0' & O"347",
    8#5447# => '0' & O"247",
    8#5450# => '0' & O"347",
    8#5451# => '0' & O"267",
    8#5452# => '0' & O"347",
    8#5453# => '0' & O"347",
    8#5454# => '0' & O"347",
    8#5455# => '0' & O"307",
    8#5456# => '0' & O"347",
    8#5457# => '0' & O"730",
    8#5460# => '1' & O"447",
    8#5461# => '0' & O"327",
    8#5462# => '0' & O"137",
    8#5463# => '0' & O"177",
    8#5464# => '0' & O"277",
    8#5465# => '1' & O"233",
    8#5466# => '0' & O"347",
    8#5467# => '0' & O"604",
    8#5470# => '1' & O"356",
    8#5471# => '0' & O"075",
    8#5472# => '1' & O"063",
    8#5473# => '0' & O"347",
    8#5474# => '0' & O"630",
    8#5475# => '1' & O"447",
    8#5476# => '0' & O"347",
    8#5477# => '0' & O"056",
    8#5500# => '0' & O"616",
    8#5501# => '0' & O"316",
    8#5502# => '0' & O"546",
    8#5503# => '1' & O"014",
    8#5504# => '0' & O"630",
    8#5505# => '0' & O"030",
    8#5506# => '0' & O"454",
    8#5507# => '0' & O"423",
    8#5510# => '0' & O"030",
    8#5511# => '1' & O"066",
    8#5512# => '0' & O"226",
    8#5513# => '0' & O"776",
    8#5514# => '1' & O"126",
    8#5515# => '0' & O"752",
    8#5516# => '1' & O"176",
    8#5517# => '0' & O"337",
    8#5520# => '1' & O"172",
    8#5521# => '1' & O"647",
    8#5522# => '1' & O"552",
    8#5523# => '1' & O"613",
    8#5524# => '1' & O"316",
    8#5525# => '1' & O"316",
    8#5526# => '1' & O"316",
    8#5527# => '1' & O"316",
    8#5530# => '1' & O"322",
    8#5531# => '1' & O"322",
    8#5532# => '0' & O"714",
    8#5533# => '0' & O"102",
    8#5534# => '0' & O"337",
    8#5535# => '0' & O"514",
    8#5536# => '0' & O"102",
    8#5537# => '0' & O"337",
    8#5540# => '0' & O"604",
    8#5541# => '1' & O"741",
    8#5542# => '1' & O"044",
    8#5543# => '0' & O"044",
    8#5544# => '0' & O"034",
    8#5545# => '1' & O"354",
    8#5546# => '0' & O"623",
    8#5547# => '0' & O"024",
    8#5550# => '1' & O"017",
    8#5551# => '1' & O"024",
    8#5552# => '0' & O"617",
    8#5553# => '0' & O"320",
    8#5554# => '1' & O"111",
    8#5555# => '0' & O"456",
    8#5556# => '0' & O"302",
    8#5557# => '1' & O"160",
    8#5560# => '1' & O"656",
    8#5561# => '1' & O"370",
    8#5562# => '1' & O"656",
    8#5563# => '1' & O"111",
    8#5564# => '1' & O"656",
    8#5565# => '1' & O"360",
    8#5566# => '1' & O"656",
    8#5567# => '0' & O"742",
    8#5570# => '0' & O"677",
    8#5571# => '0' & O"216",
    8#5572# => '0' & O"420",
    8#5573# => '1' & O"765",
    8#5574# => '1' & O"247",
    8#5575# => '0' & O"530",
    8#5576# => '1' & O"447",
    8#5577# => '0' & O"430",
    8#5600# => '1' & O"447",
    8#5601# => '0' & O"330",
    8#5602# => '1' & O"447",
    8#5603# => '1' & O"004",
    8#5604# => '1' & O"344",
    8#5605# => '1' & O"324",
    8#5606# => '0' & O"663",
    8#5607# => '0' & O"617",
    8#5610# => '0' & O"624",
    8#5611# => '0' & O"603",
    8#5612# => '0' & O"064",
    8#5613# => '0' & O"027",
    8#5614# => '1' & O"056",
    8#5615# => '0' & O"352",
    8#5616# => '1' & O"056",
    8#5617# => '0' & O"624",
    8#5620# => '0' & O"757",
    8#5621# => '0' & O"603",
    8#5622# => '1' & O"414",
    8#5623# => '1' & O"156",
    8#5624# => '1' & O"137",
    8#5625# => '1' & O"314",
    8#5626# => '0' & O"060",
    8#5627# => '1' & O"142",
    8#5630# => '1' & O"127",
    8#5631# => '0' & O"314",
    8#5632# => '0' & O"422",
    8#5633# => '0' & O"422",
    8#5634# => '0' & O"416",
    8#5635# => '0' & O"416",
    8#5636# => '1' & O"752",
    8#5637# => '1' & O"414",
    8#5640# => '0' & O"406",
    8#5641# => '1' & O"142",
    8#5642# => '1' & O"127",
    8#5643# => '1' & O"552",
    8#5644# => '1' & O"050",
    8#5645# => '1' & O"203",
    8#5646# => '1' & O"423",
    8#5647# => '1' & O"360",
    8#5650# => '1' & O"656",
    8#5651# => '0' & O"114",
    8#5652# => '1' & O"762",
    8#5653# => '1' & O"703",
    8#5654# => '0' & O"414",
    8#5655# => '1' & O"742",
    8#5656# => '0' & O"027",
    8#5657# => '0' & O"514",
    8#5660# => '1' & O"742",
    8#5661# => '0' & O"102",
    8#5662# => '1' & O"323",
    8#5663# => '0' & O"147",
    8#5664# => '1' & O"342",
    8#5665# => '0' & O"614",
    8#5666# => '1' & O"742",
    8#5667# => '0' & O"227",
    8#5670# => '0' & O"714",
    8#5671# => '1' & O"742",
    8#5672# => '0' & O"102",
    8#5673# => '1' & O"367",
    8#5674# => '0' & O"327",
    8#5675# => '1' & O"342",
    8#5676# => '1' & O"014",
    8#5677# => '1' & O"742",
    8#5700# => '1' & O"563",
    8#5701# => '1' & O"114",
    8#5702# => '1' & O"742",
    8#5703# => '1' & O"575",
    8#5704# => '0' & O"724",
    8#5705# => '1' & O"517",
    8#5706# => '1' & O"314",
    8#5707# => '0' & O"064",
    8#5710# => '0' & O"320",
    8#5711# => '1' & O"160",
    8#5712# => '1' & O"656",
    8#5713# => '0' & O"624",
    8#5714# => '1' & O"237",
    8#5715# => '1' & O"370",
    8#5716# => '1' & O"414",
    8#5717# => '0' & O"142",
    8#5720# => '0' & O"403",
    8#5721# => '1' & O"656",
    8#5722# => '0' & O"603",
    8#5723# => '0' & O"044",
    8#5724# => '0' & O"024",
    8#5725# => '1' & O"553",
    8#5726# => '1' & O"024",
    8#5727# => '1' & O"607",
    8#5730# => '0' & O"704",
    8#5731# => '0' & O"007",
    8#5732# => '1' & O"004",
    8#5733# => '1' & O"607",
    8#5734# => '1' & O"214",
    8#5735# => '0' & O"034",
    8#5736# => '1' & O"054",
    8#5737# => '1' & O"567",
    8#5740# => '0' & O"007",
    8#5741# => '1' & O"603",
    8#5742# => '0' & O"426",
    8#5743# => '1' & O"552",
    8#5744# => '0' & O"337",
    8#5745# => '0' & O"523",
    8#5746# => '1' & O"166",
    8#5747# => '1' & O"647",
    8#5750# => '0' & O"343",
    8#5751# => '1' & O"326",
    8#5752# => '1' & O"752",
    8#5753# => '1' & O"633",
    8#5754# => '0' & O"523",
    8#5755# => '1' & O"064",
    8#5756# => '0' & O"103",
    8#5757# => '0' & O"000",
    8#5760# => '1' & O"741",
    8#5761# => '0' & O"147",
    8#5762# => '0' & O"230",
    8#5763# => '1' & O"447",
    8#5764# => '0' & O"130",
    8#5765# => '1' & O"447",
    8#5766# => '0' & O"030",
    8#5767# => '1' & O"447",
    8#5770# => '1' & O"114",
    8#5771# => '1' & O"142",
    8#5772# => '1' & O"773",
    8#5773# => '1' & O"042",
    8#5774# => '0' & O"202",
    8#5775# => '0' & O"060",
    8#5776# => '0' & O"042",
    8#5777# => '1' & O"767"
  );  -- End 55 ROM

end rom_pack;

package body rom_pack is
end rom_pack;
